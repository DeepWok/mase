module llm_int #(

)(

);

scatter

matrix_mult_lp

matrix_mult_hp


gather




endmodule