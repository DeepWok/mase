`timescale 1ns / 1ps

module fixed_gqa_input_block #(
    parameter DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter DATA_IN_0_TENSOR_SIZE_DIM_1 = 20,
    parameter DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter DATA_IN_0_PARALLELISM_DIM_1 = 4,
    parameter DATA_IN_0_PRECISION_0 = 16,
    parameter DATA_IN_0_PRECISION_1 = 3,

    // Q Weights
    parameter WEIGHTS_PRE_TRANSPOSED = 0,
    parameter WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter WEIGHT_PRECISION_0 = 16,
    parameter WEIGHT_PRECISION_1 = 3,

    // K & V weights params
    localparam GROUPED_WEIGHT_TENSOR_SIZE_DIM_0 = WEIGHT_TENSOR_SIZE_DIM_0 / GROUP_SIZE,
    localparam GROUPED_WEIGHT_TENSOR_SIZE_DIM_1 = WEIGHT_TENSOR_SIZE_DIM_1,
    // Assuption: shared weights have same parallelism
    localparam GROUPED_WEIGHT_PARALLELISM_DIM_0 = WEIGHT_PARALLELISM_DIM_0,
    localparam GROUPED_WEIGHT_PARALLELISM_DIM_1 = WEIGHT_PARALLELISM_DIM_1,
    // Assuption: shared weights have same fixed point format
    localparam GROUPED_WEIGHT_PRECISION_0 = WEIGHT_PRECISION_0,
    localparam GROUPED_WEIGHT_PRECISION_1 = WEIGHT_PRECISION_1,

    parameter HAS_BIAS = 1,
    parameter BIAS_TENSOR_SIZE_DIM_0 = 64,
    parameter BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter BIAS_PARALLELISM_DIM_0 = 4,
    parameter BIAS_PARALLELISM_DIM_1 = 1,
    parameter BIAS_PRECISION_0 = 16,
    parameter BIAS_PRECISION_1 = 3,

    parameter DATA_OUT_0_TENSOR_SIZE_DIM_0 = WEIGHT_TENSOR_SIZE_DIM_0,
    parameter DATA_OUT_0_TENSOR_SIZE_DIM_1 = DATA_IN_0_TENSOR_SIZE_DIM_1,
    parameter DATA_OUT_0_PARALLELISM_DIM_0 = WEIGHT_PARALLELISM_DIM_0,
    parameter DATA_OUT_0_PARALLELISM_DIM_1 = DATA_IN_0_PARALLELISM_DIM_1,
    parameter DATA_OUT_0_PRECISION_0 = 16,
    parameter DATA_OUT_0_PRECISION_1 = 3

) (
    input logic clk,
    input logic rst,

    input logic [DATA_IN_0_PRECISION_0-1:0] data_in_0 [DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1-1:0],
    input logic data_in_0_valid,
    output logic data_in_0_ready,

    // Query weights
    input logic [WEIGHT_PRECISION_0-1:0] weight_query [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    input logic weight_query_valid,
    output logic weight_query_ready,

    // Query bias
    input logic [BIAS_PRECISION_0-1:0] bias_query [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1 -1:0],
    input logic bias_query_valid,
    output logic bias_query_ready,

    // Key weights
    input logic [WEIGHT_PRECISION_0-1:0] weight_key [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    input logic weight_key_valid,
    output logic weight_key_ready,

    // Key bias
    input logic [BIAS_PRECISION_0-1:0] bias_key [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1 -1:0],
    input logic bias_key_valid,
    output logic bias_key_ready,

    // Value weights
    input logic [WEIGHT_PRECISION_0-1:0] weight_value [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    input logic weight_value_valid,
    output logic weight_value_ready,

    // Value bias
    input logic [BIAS_PRECISION_0-1:0] bias_value [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1 -1:0],
    input logic bias_value_valid,
    output logic bias_value_ready,

    // Query
    output logic [DATA_OUT_0_PRECISION_0-1:0] data_out_query [DATA_IN_0_PARALLELISM_DIM_1 * WEIGHT_PARALLELISM_DIM_0-1:0],
    output logic data_out_query_valid,
    input logic data_out_query_ready,

    // Key
    output logic [DATA_OUT_0_PRECISION_0-1:0] data_out_key [DATA_IN_0_PARALLELISM_DIM_1 * WEIGHT_PARALLELISM_DIM_0-1:0],
    output logic data_out_key_valid,
    input logic data_out_key_ready,

    // Value
    output logic [DATA_OUT_0_PRECISION_0-1:0] data_out_value [DATA_IN_0_PARALLELISM_DIM_1 * WEIGHT_PARALLELISM_DIM_0-1:0],
    output logic data_out_value_valid,
    input logic data_out_value_ready
);

  // ! TO DO: add assertions about bias parallelism matching weight parallelism

  // * Inferred parameters
  parameter DATA_IN_0_DEPTH_DIM_1 = DATA_IN_0_TENSOR_SIZE_DIM_1 / DATA_IN_0_PARALLELISM_DIM_1;
  parameter WEIGHT_DEPTH_DIM_0 = WEIGHT_TENSOR_SIZE_DIM_0 / WEIGHT_PARALLELISM_DIM_0;

  // * Declarations
  // * =================================================================

  logic query_data_in_valid, query_data_in_ready;
  logic key_data_in_valid, key_data_in_ready;
  logic value_data_in_valid, value_data_in_ready;

  logic [DATA_OUT_0_PRECISION_0-1:0] query_buffer [DATA_IN_0_PARALLELISM_DIM_1 * WEIGHT_PARALLELISM_DIM_0-1:0];
  logic query_buffer_valid;
  logic query_buffer_ready;

  // * Instances
  // * =================================================================

  // * Split the incoming data over the QKV projections
  split_n #(
      .N(3)
  ) split_i (
      .data_in_valid (data_in_0_valid),
      .data_in_ready (data_in_0_ready),
      .data_out_valid({query_data_in_valid, key_data_in_valid, value_data_in_valid}),
      .data_out_ready({query_data_in_ready, key_data_in_ready, value_data_in_ready})
  );

  // * Query linear

//   fixed_linear #(
//       .HAS_BIAS              (HAS_BIAS),
//       .WEIGHTS_PRE_TRANSPOSED(WEIGHTS_PRE_TRANSPOSED),

//       .DATA_IN_0_PRECISION_0      (DATA_IN_0_PRECISION_0),
//       .DATA_IN_0_PRECISION_1      (DATA_IN_0_PRECISION_1),
//       .DATA_IN_0_TENSOR_SIZE_DIM_0(DATA_IN_0_TENSOR_SIZE_DIM_0),
//       .DATA_IN_0_TENSOR_SIZE_DIM_1(DATA_IN_0_TENSOR_SIZE_DIM_1),
//       .DATA_IN_0_PARALLELISM_DIM_0(DATA_IN_0_PARALLELISM_DIM_0),
//       .DATA_IN_0_PARALLELISM_DIM_1(DATA_IN_0_PARALLELISM_DIM_1),

//       .WEIGHT_PRECISION_0      (WEIGHT_PRECISION_0),
//       .WEIGHT_PRECISION_1      (WEIGHT_PRECISION_1),
//       .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
//       .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
//       .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
//       .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1),

//       .BIAS_PRECISION_0      (BIAS_PRECISION_0),
//       .BIAS_PRECISION_1      (BIAS_PRECISION_1),
//       .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
//       .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
//       .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
//       .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1),

//       .DATA_OUT_0_PRECISION_0(DATA_OUT_0_PRECISION_0),
//       .DATA_OUT_0_PRECISION_1(DATA_OUT_0_PRECISION_1)

//   ) fixed_linear_query (
//       .clk,
//       .rst,

//       // input port for data_inivations
//       .data_in_0      (data_in_0),
//       .data_in_0_valid(query_data_in_valid),
//       .data_in_0_ready(query_data_in_ready),

//       // input port for weight
//       .weight      (weight_query),
//       .weight_valid(weight_query_valid),
//       .weight_ready(weight_query_ready),

//       .bias      (bias_query),
//       .bias_valid(bias_query_valid),
//       .bias_ready(bias_query_ready),

//       .data_out_0      (query_buffer),
//       .data_out_0_valid(query_buffer_valid),
//       .data_out_0_ready(query_buffer_ready)
//   );

//   // * We must buffer the queries to latency match the key transpose path
//   // * since the matmul for QK^T buffers K^T but streams Q
//   matrix_fifo #(
//       .DATA_WIDTH(DATA_OUT_0_PRECISION_0),
//       .DIM0      (WEIGHT_PARALLELISM_DIM_0),
//       .DIM1      (DATA_IN_0_PARALLELISM_DIM_1),
//       .FIFO_SIZE (DATA_IN_0_DEPTH_DIM_1 * WEIGHT_DEPTH_DIM_0)
//   ) query_buffer_i (
//       .clk,
//       .rst,
//       .in_data  (query_buffer),
//       .in_valid (query_buffer_valid),
//       .in_ready (query_buffer_ready),
//       .out_data (data_out_query),
//       .out_valid(data_out_query_valid),
//       .out_ready(data_out_query_ready)
//   );

//   // * Key linear

//   fixed_linear #(
//       .HAS_BIAS              (HAS_BIAS),
//       .WEIGHTS_PRE_TRANSPOSED(WEIGHTS_PRE_TRANSPOSED),

//       .DATA_IN_0_PRECISION_0      (DATA_IN_0_PRECISION_0),
//       .DATA_IN_0_PRECISION_1      (DATA_IN_0_PRECISION_1),
//       .DATA_IN_0_TENSOR_SIZE_DIM_0(DATA_IN_0_TENSOR_SIZE_DIM_0),
//       .DATA_IN_0_TENSOR_SIZE_DIM_1(DATA_IN_0_TENSOR_SIZE_DIM_1),
//       .DATA_IN_0_PARALLELISM_DIM_0(DATA_IN_0_PARALLELISM_DIM_0),
//       .DATA_IN_0_PARALLELISM_DIM_1(DATA_IN_0_PARALLELISM_DIM_1),

//       .WEIGHT_PRECISION_0      (WEIGHT_PRECISION_0),
//       .WEIGHT_PRECISION_1      (WEIGHT_PRECISION_1),
//       .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
//       .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
//       .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
//       .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1),

//       .BIAS_PRECISION_0      (BIAS_PRECISION_0),
//       .BIAS_PRECISION_1      (BIAS_PRECISION_1),
//       .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
//       .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
//       .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
//       .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1),

//       .DATA_OUT_0_PRECISION_0(DATA_OUT_0_PRECISION_0),
//       .DATA_OUT_0_PRECISION_1(DATA_OUT_0_PRECISION_1)

//   ) fixed_linear_key (
//       .clk,
//       .rst,

//       // input port for data_inivations
//       .data_in_0      (data_in_0),
//       .data_in_0_valid(key_data_in_valid),
//       .data_in_0_ready(key_data_in_ready),

//       // input port for weight
//       .weight      (weight_key),
//       .weight_valid(weight_key_valid),
//       .weight_ready(weight_key_ready),

//       .bias      (bias_key),
//       .bias_valid(bias_key_valid),
//       .bias_ready(bias_key_ready),

//       .data_out_0      (data_out_key),
//       .data_out_0_valid(data_out_key_valid),
//       .data_out_0_ready(data_out_key_ready)
//   );

//   // * Value linear

//   fixed_linear #(
//       .HAS_BIAS              (HAS_BIAS),
//       .WEIGHTS_PRE_TRANSPOSED(WEIGHTS_PRE_TRANSPOSED),

//       .DATA_IN_0_PRECISION_0      (DATA_IN_0_PRECISION_0),
//       .DATA_IN_0_PRECISION_1      (DATA_IN_0_PRECISION_1),
//       .DATA_IN_0_TENSOR_SIZE_DIM_0(DATA_IN_0_TENSOR_SIZE_DIM_0),
//       .DATA_IN_0_TENSOR_SIZE_DIM_1(DATA_IN_0_TENSOR_SIZE_DIM_1),
//       .DATA_IN_0_PARALLELISM_DIM_0(DATA_IN_0_PARALLELISM_DIM_0),
//       .DATA_IN_0_PARALLELISM_DIM_1(DATA_IN_0_PARALLELISM_DIM_1),

//       .WEIGHT_PRECISION_0      (WEIGHT_PRECISION_0),
//       .WEIGHT_PRECISION_1      (WEIGHT_PRECISION_1),
//       .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
//       .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
//       .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
//       .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1),

//       .BIAS_PRECISION_0      (BIAS_PRECISION_0),
//       .BIAS_PRECISION_1      (BIAS_PRECISION_1),
//       .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
//       .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
//       .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
//       .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1),

//       .DATA_OUT_0_PRECISION_0(DATA_OUT_0_PRECISION_0),
//       .DATA_OUT_0_PRECISION_1(DATA_OUT_0_PRECISION_1)

//   ) fixed_linear_value (
//       .clk,
//       .rst,

//       // input port for data_inivations
//       .data_in_0      (data_in_0),
//       .data_in_0_valid(value_data_in_valid),
//       .data_in_0_ready(value_data_in_ready),

//       // input port for weight
//       .weight      (weight_value),
//       .weight_valid(weight_value_valid),
//       .weight_ready(weight_value_ready),

//       .bias      (bias_value),
//       .bias_valid(bias_value_valid),
//       .bias_ready(bias_value_ready),

//       .data_out_0      (data_out_value),
//       .data_out_0_valid(data_out_value_valid),
//       .data_out_0_ready(data_out_value_ready)
//   );

endmodule
