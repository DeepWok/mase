
`timescale 1ns / 1ps
/* verilator lint_off UNUSEDPARAM */
module isqrt_lut #(
    parameter DATA_IN_0_PRECISION_0  = 16,
    parameter DATA_IN_0_PRECISION_1  = 8,
    parameter DATA_OUT_0_PRECISION_0 = 16,
    parameter DATA_OUT_0_PRECISION_1 = 8
) (
    /* verilator lint_off UNUSEDSIGNAL */
    input  logic [7:0] data_in_0,
    output logic [7:0] data_out_0
);

  always_comb begin
    case (data_in_0)
      8'b00000000: data_out_0 = 8'b01111111;
      8'b00000001: data_out_0 = 8'b01111111;
      8'b00000010: data_out_0 = 8'b01111111;
      8'b00000011: data_out_0 = 8'b01111111;
      8'b00000100: data_out_0 = 8'b01111111;
      8'b00000101: data_out_0 = 8'b01111111;
      8'b00000110: data_out_0 = 8'b01111111;
      8'b00000111: data_out_0 = 8'b01111111;
      8'b00001000: data_out_0 = 8'b01111111;
      8'b00001001: data_out_0 = 8'b01111000;
      8'b00001010: data_out_0 = 8'b01110010;
      8'b00001011: data_out_0 = 8'b01101101;
      8'b00001100: data_out_0 = 8'b01101000;
      8'b00001101: data_out_0 = 8'b01100100;
      8'b00001110: data_out_0 = 8'b01100000;
      8'b00001111: data_out_0 = 8'b01011101;
      8'b00010000: data_out_0 = 8'b01011010;
      8'b00010001: data_out_0 = 8'b01010111;
      8'b00010010: data_out_0 = 8'b01010101;
      8'b00010011: data_out_0 = 8'b01010011;
      8'b00010100: data_out_0 = 8'b01010000;
      8'b00010101: data_out_0 = 8'b01001111;
      8'b00010110: data_out_0 = 8'b01001101;
      8'b00010111: data_out_0 = 8'b01001011;
      8'b00011000: data_out_0 = 8'b01001001;
      8'b00011001: data_out_0 = 8'b01001000;
      8'b00011010: data_out_0 = 8'b01000111;
      8'b00011011: data_out_0 = 8'b01000101;
      8'b00011100: data_out_0 = 8'b01000100;
      8'b00011101: data_out_0 = 8'b01000011;
      8'b00011110: data_out_0 = 8'b01000010;
      8'b00011111: data_out_0 = 8'b01000001;
      8'b00100000: data_out_0 = 8'b00111111;
      8'b00100001: data_out_0 = 8'b00111111;
      8'b00100010: data_out_0 = 8'b00111110;
      8'b00100011: data_out_0 = 8'b00111101;
      8'b00100100: data_out_0 = 8'b00111100;
      8'b00100101: data_out_0 = 8'b00111011;
      8'b00100110: data_out_0 = 8'b00111010;
      8'b00100111: data_out_0 = 8'b00111001;
      8'b00101000: data_out_0 = 8'b00111001;
      8'b00101001: data_out_0 = 8'b00111000;
      8'b00101010: data_out_0 = 8'b00110111;
      8'b00101011: data_out_0 = 8'b00110111;
      8'b00101100: data_out_0 = 8'b00110110;
      8'b00101101: data_out_0 = 8'b00110101;
      8'b00101110: data_out_0 = 8'b00110101;
      8'b00101111: data_out_0 = 8'b00110100;
      8'b00110000: data_out_0 = 8'b00110100;
      8'b00110001: data_out_0 = 8'b00110011;
      8'b00110010: data_out_0 = 8'b00110011;
      8'b00110011: data_out_0 = 8'b00110010;
      8'b00110100: data_out_0 = 8'b00110010;
      8'b00110101: data_out_0 = 8'b00110001;
      8'b00110110: data_out_0 = 8'b00110001;
      8'b00110111: data_out_0 = 8'b00110000;
      8'b00111000: data_out_0 = 8'b00110000;
      8'b00111001: data_out_0 = 8'b00101111;
      8'b00111010: data_out_0 = 8'b00101111;
      8'b00111011: data_out_0 = 8'b00101111;
      8'b00111100: data_out_0 = 8'b00101110;
      8'b00111101: data_out_0 = 8'b00101110;
      8'b00111110: data_out_0 = 8'b00101101;
      8'b00111111: data_out_0 = 8'b00101101;
      8'b01000000: data_out_0 = 8'b00101101;
      8'b01000001: data_out_0 = 8'b00101100;
      8'b01000010: data_out_0 = 8'b00101100;
      8'b01000011: data_out_0 = 8'b00101100;
      8'b01000100: data_out_0 = 8'b00101011;
      8'b01000101: data_out_0 = 8'b00101011;
      8'b01000110: data_out_0 = 8'b00101011;
      8'b01000111: data_out_0 = 8'b00101010;
      8'b01001000: data_out_0 = 8'b00101010;
      8'b01001001: data_out_0 = 8'b00101010;
      8'b01001010: data_out_0 = 8'b00101010;
      8'b01001011: data_out_0 = 8'b00101001;
      8'b01001100: data_out_0 = 8'b00101001;
      8'b01001101: data_out_0 = 8'b00101001;
      8'b01001110: data_out_0 = 8'b00101000;
      8'b01001111: data_out_0 = 8'b00101000;
      8'b01010000: data_out_0 = 8'b00101000;
      8'b01010001: data_out_0 = 8'b00101000;
      8'b01010010: data_out_0 = 8'b00100111;
      8'b01010011: data_out_0 = 8'b00100111;
      8'b01010100: data_out_0 = 8'b00100111;
      8'b01010101: data_out_0 = 8'b00100111;
      8'b01010110: data_out_0 = 8'b00100111;
      8'b01010111: data_out_0 = 8'b00100110;
      8'b01011000: data_out_0 = 8'b00100110;
      8'b01011001: data_out_0 = 8'b00100110;
      8'b01011010: data_out_0 = 8'b00100110;
      8'b01011011: data_out_0 = 8'b00100101;
      8'b01011100: data_out_0 = 8'b00100101;
      8'b01011101: data_out_0 = 8'b00100101;
      8'b01011110: data_out_0 = 8'b00100101;
      8'b01011111: data_out_0 = 8'b00100101;
      8'b01100000: data_out_0 = 8'b00100100;
      8'b01100001: data_out_0 = 8'b00100100;
      8'b01100010: data_out_0 = 8'b00100100;
      8'b01100011: data_out_0 = 8'b00100100;
      8'b01100100: data_out_0 = 8'b00100100;
      8'b01100101: data_out_0 = 8'b00100100;
      8'b01100110: data_out_0 = 8'b00100011;
      8'b01100111: data_out_0 = 8'b00100011;
      8'b01101000: data_out_0 = 8'b00100011;
      8'b01101001: data_out_0 = 8'b00100011;
      8'b01101010: data_out_0 = 8'b00100011;
      8'b01101011: data_out_0 = 8'b00100010;
      8'b01101100: data_out_0 = 8'b00100010;
      8'b01101101: data_out_0 = 8'b00100010;
      8'b01101110: data_out_0 = 8'b00100010;
      8'b01101111: data_out_0 = 8'b00100010;
      8'b01110000: data_out_0 = 8'b00100010;
      8'b01110001: data_out_0 = 8'b00100010;
      8'b01110010: data_out_0 = 8'b00100001;
      8'b01110011: data_out_0 = 8'b00100001;
      8'b01110100: data_out_0 = 8'b00100001;
      8'b01110101: data_out_0 = 8'b00100001;
      8'b01110110: data_out_0 = 8'b00100001;
      8'b01110111: data_out_0 = 8'b00100001;
      8'b01111000: data_out_0 = 8'b00100001;
      8'b01111001: data_out_0 = 8'b00100000;
      8'b01111010: data_out_0 = 8'b00100000;
      8'b01111011: data_out_0 = 8'b00100000;
      8'b01111100: data_out_0 = 8'b00100000;
      8'b01111101: data_out_0 = 8'b00100000;
      8'b01111110: data_out_0 = 8'b00100000;
      8'b01111111: data_out_0 = 8'b00100000;
      default: data_out_0 = 8'b0;
    endcase
  end
endmodule
