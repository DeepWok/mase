// File: mxint_vit_attention.sv
module mxint_vit_attention_wrap #(
    parameter DATA_IN_0_PRECISION_0 = 8,
    parameter DATA_IN_0_PRECISION_1 = 8,
    parameter DATA_IN_0_TENSOR_SIZE_DIM_0 = 12,
    parameter DATA_IN_0_PARALLELISM_DIM_0 = 2,
    parameter DATA_IN_0_TENSOR_SIZE_DIM_1 = 10,
    parameter DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter DATA_IN_0_TENSOR_SIZE_DIM_2 = 1,
    parameter DATA_IN_0_PARALLELISM_DIM_2 = 1,
    parameter QUERY_WEIGHT_PRECISION_0 = 8,
    parameter QUERY_WEIGHT_PRECISION_1 = 4,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 12,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = 2,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 12,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = 2,
    parameter QUERY_BIAS_PRECISION_0 = 4,
    parameter QUERY_BIAS_PRECISION_1 = 8,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0 = 12,
    parameter QUERY_BIAS_PARALLELISM_DIM_0 = 2,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter KEY_WEIGHT_PRECISION_0 = 8,
    parameter KEY_WEIGHT_PRECISION_1 = 4,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 12,
    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = 2,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 12,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = 2,
    parameter KEY_BIAS_PRECISION_0 = 4,
    parameter KEY_BIAS_PRECISION_1 = 8,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0 = 12,
    parameter KEY_BIAS_PARALLELISM_DIM_0 = 2,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter VALUE_WEIGHT_PRECISION_0 = 8,
    parameter VALUE_WEIGHT_PRECISION_1 = 4,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 12,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = 2,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 12,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = 2,
    parameter VALUE_BIAS_PRECISION_0 = 4,
    parameter VALUE_BIAS_PRECISION_1 = 8,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0 = 12,
    parameter VALUE_BIAS_PARALLELISM_DIM_0 = 2,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter PROJ_WEIGHT_PRECISION_0 = 8,
    parameter PROJ_WEIGHT_PRECISION_1 = 4,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 12,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = 2,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 12,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = 2,
    parameter PROJ_BIAS_PRECISION_0 = 4,
    parameter PROJ_BIAS_PRECISION_1 = 8,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0 = 12,
    parameter PROJ_BIAS_PARALLELISM_DIM_0 = 2,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter DATA_OUT_0_PRECISION_0 = 4,
    parameter DATA_OUT_0_PRECISION_1 = 8,
    parameter DATA_OUT_0_TENSOR_SIZE_DIM_0 = 12,
    parameter DATA_OUT_0_PARALLELISM_DIM_0 = 2,
    parameter DATA_OUT_0_TENSOR_SIZE_DIM_1 = 10,
    parameter DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter DATA_OUT_0_TENSOR_SIZE_DIM_2 = 1,
    parameter DATA_OUT_0_PARALLELISM_DIM_2 = 1,
    parameter NUM_HEADS = 3,
    parameter HAS_BIAS = 1,
    localparam WEIGHT_PRECISION_0 = QUERY_WEIGHT_PRECISION_0,
    localparam WEIGHT_PRECISION_1 = QUERY_WEIGHT_PRECISION_1,
    localparam BIAS_PRECISION_0 = QUERY_BIAS_PRECISION_0,
    localparam BIAS_PRECISION_1 = QUERY_BIAS_PRECISION_1,
    localparam WEIGHT_PROJ_PRECISION_0 = PROJ_WEIGHT_PRECISION_0,
    localparam WEIGHT_PROJ_PRECISION_1 = PROJ_WEIGHT_PRECISION_1,
    localparam BIAS_PROJ_PRECISION_0 = PROJ_BIAS_PRECISION_0,
    localparam BIAS_PROJ_PRECISION_1 = PROJ_BIAS_PRECISION_1,
    localparam WEIGHT_TENSOR_SIZE_DIM_0 = QUERY_WEIGHT_TENSOR_SIZE_DIM_0,
    localparam WEIGHT_TENSOR_SIZE_DIM_1 = QUERY_WEIGHT_TENSOR_SIZE_DIM_1,
    localparam WEIGHT_PARALLELISM_DIM_0 = QUERY_WEIGHT_PARALLELISM_DIM_0,
    localparam WEIGHT_PARALLELISM_DIM_1 = QUERY_WEIGHT_PARALLELISM_DIM_1,
    localparam BIAS_TENSOR_SIZE_DIM_0 = QUERY_BIAS_TENSOR_SIZE_DIM_0,
    localparam BIAS_TENSOR_SIZE_DIM_1 = QUERY_BIAS_TENSOR_SIZE_DIM_1,
    localparam BIAS_PARALLELISM_DIM_0 = QUERY_BIAS_PARALLELISM_DIM_0,
    localparam BIAS_PARALLELISM_DIM_1 = QUERY_BIAS_PARALLELISM_DIM_1,
    localparam WEIGHT_PROJ_TENSOR_SIZE_DIM_0 = PROJ_WEIGHT_TENSOR_SIZE_DIM_0,
    localparam WEIGHT_PROJ_TENSOR_SIZE_DIM_1 = PROJ_WEIGHT_TENSOR_SIZE_DIM_1,
    localparam WEIGHT_PROJ_PARALLELISM_DIM_0 = PROJ_WEIGHT_PARALLELISM_DIM_0,
    localparam WEIGHT_PROJ_PARALLELISM_DIM_1 = PROJ_WEIGHT_PARALLELISM_DIM_1,
    localparam BIAS_PROJ_TENSOR_SIZE_DIM_0 = PROJ_BIAS_TENSOR_SIZE_DIM_0,
    localparam BIAS_PROJ_TENSOR_SIZE_DIM_1 = PROJ_BIAS_TENSOR_SIZE_DIM_1,
    localparam BIAS_PROJ_PARALLELISM_DIM_0 = PROJ_BIAS_PARALLELISM_DIM_0,
    localparam BIAS_PROJ_PARALLELISM_DIM_1 = PROJ_BIAS_PARALLELISM_DIM_1,
    localparam QKV_PRECISION_0 = DATA_IN_0_PRECISION_0,
    localparam QKV_PRECISION_1 = DATA_IN_0_PRECISION_1
) (
    input logic clk,
    input logic rst,

    input logic [DATA_IN_0_PRECISION_0-1:0] mdata_in_0 [DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1-1:0],
    input logic [DATA_IN_0_PRECISION_1-1:0] edata_in_0,
    input logic data_in_0_valid,
    output logic data_in_0_ready,

    // Query weights
    input logic [WEIGHT_PRECISION_0-1:0] mquery_weight [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    input logic [WEIGHT_PRECISION_1-1:0] equery_weight,
    input logic query_weight_valid,
    output logic query_weight_ready,

    // Query bias
    input logic [BIAS_PRECISION_0-1:0] mquery_bias [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1 -1:0],
    input logic [BIAS_PRECISION_1-1:0] equery_bias,
    input logic query_bias_valid,
    output logic query_bias_ready,

    // Key weights
    input logic [WEIGHT_PRECISION_0-1:0] mkey_weight [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    input logic [WEIGHT_PRECISION_1-1:0] ekey_weight,
    input logic key_weight_valid,
    output logic key_weight_ready,

    // Key bias
    input logic [BIAS_PRECISION_0-1:0] mkey_bias [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1 -1:0],
    input logic [BIAS_PRECISION_1-1:0] ekey_bias,
    input logic key_bias_valid,
    output logic key_bias_ready,

    // Value weights
    input logic [WEIGHT_PRECISION_0-1:0] mvalue_weight [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    input logic [WEIGHT_PRECISION_1-1:0] evalue_weight,
    input logic value_weight_valid,
    output logic value_weight_ready,

    // Value bias
    input logic [BIAS_PRECISION_0-1:0] mvalue_bias [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1 -1:0],
    input logic [BIAS_PRECISION_1-1:0] evalue_bias,
    input logic value_bias_valid,
    output logic value_bias_ready,

    // Proj weights
    input logic [WEIGHT_PROJ_PRECISION_0-1:0] mproj_weight [WEIGHT_PROJ_PARALLELISM_DIM_0 * WEIGHT_PROJ_PARALLELISM_DIM_1-1:0],
    input logic [WEIGHT_PROJ_PRECISION_1-1:0] eproj_weight,
    input logic proj_weight_valid,
    output logic proj_weight_ready,

    // Proj bias
    input logic [BIAS_PROJ_PRECISION_0-1:0] mproj_bias [BIAS_PROJ_PARALLELISM_DIM_0 * BIAS_PROJ_PARALLELISM_DIM_1 -1:0],
    input logic [BIAS_PROJ_PRECISION_1-1:0] eproj_bias,
    input logic proj_bias_valid,
    output logic proj_bias_ready,

    output logic [DATA_OUT_0_PRECISION_0-1:0] mdata_out_0 [DATA_OUT_0_PARALLELISM_DIM_0*DATA_OUT_0_PARALLELISM_DIM_1-1:0],
    output logic [DATA_OUT_0_PRECISION_1-1:0] edata_out_0,
    output logic data_out_0_valid,
    input logic data_out_0_ready
);
    // Internal logic here (if any)
        mxint_vit_attention #(
        .NUM_HEADS(NUM_HEADS),
        .DATA_IN_0_TENSOR_SIZE_DIM_0(DATA_IN_0_TENSOR_SIZE_DIM_0),
        .DATA_IN_0_TENSOR_SIZE_DIM_1(DATA_IN_0_TENSOR_SIZE_DIM_1),
        .DATA_IN_0_PARALLELISM_DIM_0(DATA_IN_0_PARALLELISM_DIM_0),
        .DATA_IN_0_PARALLELISM_DIM_1(DATA_IN_0_PARALLELISM_DIM_1),
        .DATA_IN_0_PRECISION_0(DATA_IN_0_PRECISION_0),
        .DATA_IN_0_PRECISION_1(DATA_IN_0_PRECISION_1),
        .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
        .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
        .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
        .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1),
        .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
        .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
        .HAS_BIAS(HAS_BIAS),
        .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
        .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
        .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
        .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1),
        .BIAS_PRECISION_0(BIAS_PRECISION_0),
        .BIAS_PRECISION_1(BIAS_PRECISION_1),
        .QKV_PRECISION_0(QKV_PRECISION_0),
        .QKV_PRECISION_1(QKV_PRECISION_1),
        .WEIGHT_PROJ_PRECISION_0(WEIGHT_PROJ_PRECISION_0),
        .WEIGHT_PROJ_PRECISION_1(WEIGHT_PROJ_PRECISION_1),
        .BIAS_PROJ_PRECISION_0(BIAS_PROJ_PRECISION_0),
        .BIAS_PROJ_PRECISION_1(BIAS_PROJ_PRECISION_1),
        .WEIGHT_PROJ_TENSOR_SIZE_DIM_0(WEIGHT_PROJ_TENSOR_SIZE_DIM_0),
        .WEIGHT_PROJ_TENSOR_SIZE_DIM_1(WEIGHT_PROJ_TENSOR_SIZE_DIM_1),
        .WEIGHT_PROJ_PARALLELISM_DIM_0(WEIGHT_PROJ_PARALLELISM_DIM_0),
        .WEIGHT_PROJ_PARALLELISM_DIM_1(WEIGHT_PROJ_PARALLELISM_DIM_1),
        .BIAS_PROJ_TENSOR_SIZE_DIM_0(BIAS_PROJ_TENSOR_SIZE_DIM_0),
        .BIAS_PROJ_TENSOR_SIZE_DIM_1(BIAS_PROJ_TENSOR_SIZE_DIM_1),
        .BIAS_PROJ_PARALLELISM_DIM_0(BIAS_PROJ_PARALLELISM_DIM_0),
        .BIAS_PROJ_PARALLELISM_DIM_1(BIAS_PROJ_PARALLELISM_DIM_1),
        .DATA_OUT_0_TENSOR_SIZE_DIM_0(DATA_OUT_0_TENSOR_SIZE_DIM_0),
        .DATA_OUT_0_TENSOR_SIZE_DIM_1(DATA_OUT_0_TENSOR_SIZE_DIM_1),
        .DATA_OUT_0_PARALLELISM_DIM_0(DATA_OUT_0_PARALLELISM_DIM_0),
        .DATA_OUT_0_PARALLELISM_DIM_1(DATA_OUT_0_PARALLELISM_DIM_1),
        .DATA_OUT_0_PRECISION_0(DATA_OUT_0_PRECISION_0),
        .DATA_OUT_0_PRECISION_1(DATA_OUT_0_PRECISION_1)
    ) mxint_vit_attention_inst (
        .clk(clk),
        .rst(rst),
        .mdata_in_0(mdata_in_0),
        .edata_in_0(edata_in_0),
        .data_in_0_valid(data_in_0_valid),
        .data_in_0_ready(data_in_0_ready),

        // Query weights
        .mweight_query(mquery_weight),
        .eweight_query(equery_weight),
        .query_weight_valid(query_weight_valid),
        .query_weight_ready(query_weight_ready),

        // Query bias
        .mquery_bias(mquery_bias),
        .equery_bias(equery_bias),
        .query_bias_valid(query_bias_valid),
        .query_bias_ready(query_bias_ready),

        // Key weights
        .mkey_weight(mkey_weight),
        .ekey_weight(ekey_weight),
        .key_weight_valid(key_weight_valid),
        .key_weight_ready(key_weight_ready),

        // Key bias
        .mkey_bias(mkey_bias),
        .ekey_bias(ekey_bias),
        .key_bias_valid(key_bias_valid),
        .key_bias_ready(key_bias_ready),

        // Value weights
        .mvalue_weight(mvalue_weight),
        .evalue_weight(evalue_weight),
        .value_weight_valid(value_weight_valid),
        .value_weight_ready(value_weight_ready),

        // Value bias
        .mvalue_bias(mvalue_bias),
        .evalue_bias(evalue_bias),
        .value_bias_valid(value_bias_valid),
        .value_bias_ready(value_bias_ready),

        // Proj weights
        .mproj_weight(mproj_weight),
        .eproj_weight(eproj_weight),
        .proj_weight_valid(proj_weight_valid),
        .proj_weight_ready(proj_weight_ready),

        // Proj bias
        .mproj_bias(mproj_bias),
        .eproj_bias(eproj_bias),
        .proj_bias_valid(proj_bias_valid),
        .proj_bias_ready(proj_bias_ready),

        .mdata_out_0(mdata_out_0),
        .edata_out_0(edata_out_0),
        .data_out_0_valid(data_out_0_valid),
        .data_out_0_ready(data_out_0_ready)
    );

endmodule