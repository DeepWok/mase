
    
`timescale 1ns/1ps
module top #(
    parameter REPEAT_TIMES = 1,
    parameter fork2_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_0_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_0_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_0_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_1_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_1_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_1_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_1_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_1_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_1_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_1_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_1_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_0_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_0_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_0_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_0_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_2_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_2_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_2_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_2_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_2_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_2_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_2_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_2_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_2_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_2_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_1_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_1_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_1_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_3_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_3_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_3_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_3_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_3_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_3_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_3_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_3_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_3_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_3_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_3_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_3_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_3_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_3_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_3_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_3_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_3_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_3_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_1_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_1_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_1_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_1_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_4_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_4_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_4_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_4_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_4_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_4_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_4_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_4_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_4_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_4_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_4_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_4_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_4_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_4_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_4_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_4_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_4_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_4_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_2_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_2_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_2_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_5_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_5_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_5_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_5_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_5_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_5_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_5_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_5_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_5_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_5_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_5_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_5_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_5_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_5_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_5_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_5_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_5_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_5_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_2_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_2_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_2_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_2_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_6_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_6_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_6_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_6_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_6_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_6_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_6_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_6_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_6_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_6_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_6_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_6_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_6_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_6_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_6_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_6_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_6_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_6_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_3_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_3_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_3_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_7_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_7_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_7_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_7_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_7_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_7_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_7_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_7_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_7_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_7_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_7_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_7_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_7_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_7_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_7_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_7_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_7_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_7_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_3_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_3_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_3_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_3_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_8_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_8_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_8_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_8_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_8_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_8_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_8_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_8_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_8_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_8_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_8_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_8_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_8_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_8_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_8_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_8_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_8_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_8_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_4_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_4_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_4_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_9_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_9_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_9_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_9_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_9_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_9_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_9_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_9_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_9_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_9_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_9_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_9_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_9_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_9_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_9_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_9_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_9_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_9_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_4_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_4_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_4_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_4_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_10_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_10_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_10_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_10_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_10_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_10_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_10_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_10_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_10_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_10_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_10_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_10_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_10_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_10_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_10_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_10_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_10_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_10_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_5_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_5_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_5_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_11_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_11_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_11_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_11_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_11_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_11_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_11_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_11_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_11_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_11_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_11_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_11_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_11_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_11_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_11_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_11_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_11_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_11_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_5_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_5_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_5_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_5_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_12_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_12_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_12_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_12_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_12_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_12_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_12_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_12_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_12_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_12_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_12_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_12_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_12_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_12_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_12_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_12_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_12_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_12_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_6_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_6_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_6_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_13_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_13_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_13_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_13_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_13_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_13_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_13_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_13_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_13_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_13_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_13_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_13_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_13_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_13_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_13_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_13_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_13_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_13_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_6_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_6_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_6_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_6_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_14_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_14_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_14_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_14_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_14_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_14_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_14_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_14_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_14_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_14_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_14_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_14_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_14_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_14_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_14_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_14_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_14_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_14_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_7_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_7_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_7_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_15_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_15_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_15_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_15_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_15_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_15_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_15_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_15_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_15_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_15_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_15_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_15_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_15_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_15_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_15_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_15_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_15_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_15_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_7_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_7_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_7_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_7_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_16_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_16_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_16_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_16_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_16_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_16_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_16_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_16_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_16_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_16_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_16_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_16_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_16_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_16_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_16_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_16_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_16_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_16_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_8_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_8_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_8_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_17_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_17_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_17_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_17_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_17_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_17_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_17_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_17_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_17_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_17_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_17_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_17_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_17_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_17_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_17_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_17_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_17_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_17_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_8_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_8_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_8_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_8_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_18_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_18_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_18_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_18_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_18_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_18_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_18_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_18_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_18_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_18_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_18_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_18_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_18_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_18_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_18_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_18_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_18_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_18_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_9_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_9_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_9_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_19_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_19_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_19_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_19_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_19_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_19_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_19_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_19_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_19_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_19_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_19_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_19_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_19_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_19_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_19_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_19_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_19_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_19_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_9_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_9_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_9_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_9_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_20_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_20_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_20_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_20_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_20_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_20_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_20_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_20_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_20_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_20_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_20_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_20_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_20_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_20_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_20_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_20_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_20_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_20_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_10_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_10_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_10_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_21_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_21_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_21_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_21_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_21_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_21_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_21_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_21_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_21_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_21_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_21_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_21_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_21_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_21_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_21_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_21_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_21_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_21_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_10_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_10_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_10_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_10_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_22_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_22_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_22_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_22_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_22_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_22_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_22_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_22_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_22_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_22_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_22_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_22_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_22_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_22_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_22_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_22_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_22_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_22_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_linear1_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter folded_blocks_0_stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_linear2_WEIGHT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter folded_blocks_0_stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_BIAS_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_norm1_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_norm1_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm1_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_11_norm1_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm1_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_11_norm1_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_11_norm1_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_23_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_23_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_23_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_23_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_23_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_23_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_23_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_23_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_23_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_23_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_23_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_23_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_23_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_23_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_23_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_23_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_23_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_23_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_WEIGHT_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_norm2_WEIGHT_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_BIAS_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_norm2_BIAS_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_ELEMENTWISE_AFFINE = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_HAS_BIAS = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_norm2_ISQRT_IN_PRECISION_0 = 8,
    parameter folded_blocks_0_stream_blocks_11_norm2_ISQRT_IN_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_norm2_ISQRT_OUT_PRECISION_0 = 16,
    parameter folded_blocks_0_stream_blocks_11_norm2_ISQRT_OUT_PRECISION_1 = 8,
    parameter folded_blocks_0_stream_blocks_11_norm2_ISQRT_OUT_EXPONENT_PRECISION_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter folded_blocks_0_stream_blocks_11_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter DATA_IN_0_PRECISION_0 = 6,
    parameter DATA_IN_0_PRECISION_1 = 4,
    parameter DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter DATA_OUT_0_PRECISION_0 = 6,
    parameter DATA_OUT_0_PRECISION_1 = 4,
    parameter DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter DATA_OUT_0_PARALLELISM_DIM_1 = 1
) (
    input clk,
    input rst,
    input logic [DATA_IN_0_PRECISION_0-1:0]  mdata_in_0       [DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1-1:0],
    input logic [DATA_IN_0_PRECISION_1-1:0]  edata_in_0,
    input logic                             data_in_0_valid,
    output logic                             data_in_0_ready,
    output logic [DATA_IN_0_PRECISION_0-1:0]  mdata_out_0       [DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1-1:0],
    output logic [DATA_IN_0_PRECISION_1-1:0]  edata_out_0,
    output logic                             data_out_0_valid,
    input logic                             data_out_0_ready
);
localparam IMAGE_DEPTH = DATA_IN_0_TENSOR_SIZE_DIM_0 * DATA_IN_0_TENSOR_SIZE_DIM_1 / (DATA_IN_0_PARALLELISM_DIM_1*DATA_IN_0_PARALLELISM_DIM_0);
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
localparam MAN_WIDTH = DATA_IN_0_PRECISION_0;
localparam EXP_WIDTH = DATA_IN_0_PRECISION_1;
localparam IN_SIZE = DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1;


logic [DATA_IN_0_PRECISION_0-1:0]  top_block_mdata_in_0       [DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [DATA_IN_0_PRECISION_1-1:0]  top_block_edata_in_0;
logic                             top_block_data_in_0_valid;
logic                             top_block_data_in_0_ready;

logic [DATA_IN_0_PRECISION_0-1:0]  top_block_mdata_out_0       [DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [DATA_IN_0_PRECISION_1-1:0]  top_block_edata_out_0;
logic                             top_block_data_out_0_valid;
logic                             top_block_data_out_0_ready;

logic [DATA_IN_0_PRECISION_0-1:0]  a_fifo_mdata_out_0       [DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [DATA_IN_0_PRECISION_1-1:0]  a_fifo_edata_out_0;
logic                             a_fifo_data_out_0_valid;
logic                             a_fifo_data_out_0_ready;

logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter_in, counter_out;
always_ff @(posedge clk)
    if (rst) counter_in <= 0;
    else
        if (counter_in == COUNTER_DEPTH) counter_in <= 0;
        else if (top_block_data_in_0_valid && top_block_data_in_0_ready) counter_in <= counter_in + 1;

always_ff @(posedge clk)
    if (rst) counter_out <= 0;
    else
        if (counter_out == COUNTER_DEPTH) counter_out <= 0;
        else if (a_fifo_data_out_0_valid && a_fifo_data_out_0_ready) counter_out <= counter_out + 1;

top_block top_block_inst (
    .clk(clk),
    .rst(rst),
    .mdata_in_0(top_block_mdata_in_0),
    .edata_in_0(top_block_edata_in_0),
    .data_in_0_valid(top_block_data_in_0_valid),
    .data_in_0_ready(top_block_data_in_0_ready),
    .mdata_out_0(top_block_mdata_out_0),
    .edata_out_0(top_block_edata_out_0),
    .data_out_0_valid(top_block_data_out_0_valid),
    .data_out_0_ready(top_block_data_out_0_ready)
);


  unpacked_mx_fifo #(
    .MAN_WIDTH(DATA_IN_0_PRECISION_0),
    .EXP_WIDTH(DATA_IN_0_PRECISION_1), 
    .IN_SIZE(DATA_IN_0_PARALLELISM_DIM_0 * DATA_IN_0_PARALLELISM_DIM_1),
    .DEPTH(IMAGE_DEPTH)  // Minimum depth for breaking timing path
  ) data_fifo (
    .clk(clk),
    .rst(rst),
    .mdata_in(top_block_mdata_out_0),
    .edata_in(top_block_edata_out_0),
    .data_in_valid(top_block_data_out_0_valid),
    .data_in_ready(top_block_data_out_0_ready),
    .mdata_out(a_fifo_mdata_out_0),
    .edata_out(a_fifo_edata_out_0),
    .data_out_valid(a_fifo_data_out_0_valid),
    .data_out_ready(a_fifo_data_out_0_ready)
  );

always_comb begin
    top_block_mdata_in_0 = (counter_in < IMAGE_DEPTH)? mdata_in_0: a_fifo_mdata_out_0;
    top_block_edata_in_0 = (counter_in < IMAGE_DEPTH)? edata_in_0: a_fifo_edata_out_0;
    top_block_data_in_0_valid = (counter_in < IMAGE_DEPTH)? data_in_0_valid: a_fifo_data_out_0_valid;
    data_in_0_ready = (counter_in < IMAGE_DEPTH)? top_block_data_in_0_ready: 1'b0;
end
always_comb begin
    mdata_out_0 = a_fifo_mdata_out_0;
    edata_out_0 = a_fifo_edata_out_0;
    data_out_0_valid = (counter_out < (REPEAT_TIMES - 1)*IMAGE_DEPTH)? 0: a_fifo_data_out_0_valid;
    a_fifo_data_out_0_ready = (counter_out >= (REPEAT_TIMES - 1)*IMAGE_DEPTH)? data_out_0_ready: (counter_in < IMAGE_DEPTH) ? 0 : top_block_data_in_0_ready; 
end
endmodule
    
    
// =====================================
//     Mase Hardware
//     Model: top_block
//     09/01/2025 01:34:32
// =====================================
`timescale 1ns/1ps
module top_block #(
    parameter fork2_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_0_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_0_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_0_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_0_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_0_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_0_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_0_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_0_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_0_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_0_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_0_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_0_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_0_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_0_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_0_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_0_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_0_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_0_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_0_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_0_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_0_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_0_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_0_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_0_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_0_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_0_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_0_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_0_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_0_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_0_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_0_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_0_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_0_norm1_HAS_BIAS = 1,
    parameter stream_blocks_0_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_0_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_0_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_0_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_0_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_0_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_0_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_0_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_0_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_1_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_1_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_1_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_1_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_1_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_1_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_1_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_1_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_0_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_0_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_0_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_0_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_0_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_0_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_0_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_0_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_0_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_0_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_0_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_0_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_0_norm2_HAS_BIAS = 1,
    parameter stream_blocks_0_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_0_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_0_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_0_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_0_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_0_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_0_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_0_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_0_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_0_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_0_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_0_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_0_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_2_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_2_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_2_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_2_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_2_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_2_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_2_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_2_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_2_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_2_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_1_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_1_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_1_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_1_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_1_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_1_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_1_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_1_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_1_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_1_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_1_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_1_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_1_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_1_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_1_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_1_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_1_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_1_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_1_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_1_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_1_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_1_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_1_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_1_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_1_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_1_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_1_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_1_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_1_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_1_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_1_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_1_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_1_norm1_HAS_BIAS = 1,
    parameter stream_blocks_1_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_1_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_1_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_1_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_1_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_1_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_1_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_1_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_1_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_3_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_3_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_3_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_3_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_3_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_3_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_3_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_3_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_3_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_3_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_3_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_3_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_3_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_3_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_3_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_3_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_3_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_3_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_1_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_1_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_1_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_1_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_1_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_1_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_1_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_1_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_1_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_1_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_1_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_1_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_1_norm2_HAS_BIAS = 1,
    parameter stream_blocks_1_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_1_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_1_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_1_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_1_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_1_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_1_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_1_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_1_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_1_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_1_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_1_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_1_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_4_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_4_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_4_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_4_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_4_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_4_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_4_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_4_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_4_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_4_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_4_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_4_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_4_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_4_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_4_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_4_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_4_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_4_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_2_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_2_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_2_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_2_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_2_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_2_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_2_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_2_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_2_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_2_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_2_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_2_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_2_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_2_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_2_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_2_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_2_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_2_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_2_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_2_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_2_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_2_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_2_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_2_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_2_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_2_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_2_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_2_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_2_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_2_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_2_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_2_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_2_norm1_HAS_BIAS = 1,
    parameter stream_blocks_2_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_2_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_2_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_2_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_2_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_2_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_2_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_2_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_2_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_5_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_5_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_5_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_5_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_5_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_5_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_5_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_5_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_5_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_5_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_5_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_5_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_5_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_5_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_5_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_5_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_5_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_5_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_2_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_2_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_2_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_2_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_2_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_2_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_2_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_2_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_2_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_2_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_2_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_2_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_2_norm2_HAS_BIAS = 1,
    parameter stream_blocks_2_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_2_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_2_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_2_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_2_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_2_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_2_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_2_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_2_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_2_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_2_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_2_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_2_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_6_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_6_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_6_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_6_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_6_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_6_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_6_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_6_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_6_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_6_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_6_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_6_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_6_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_6_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_6_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_6_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_6_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_6_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_3_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_3_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_3_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_3_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_3_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_3_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_3_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_3_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_3_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_3_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_3_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_3_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_3_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_3_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_3_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_3_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_3_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_3_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_3_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_3_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_3_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_3_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_3_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_3_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_3_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_3_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_3_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_3_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_3_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_3_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_3_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_3_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_3_norm1_HAS_BIAS = 1,
    parameter stream_blocks_3_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_3_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_3_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_3_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_3_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_3_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_3_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_3_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_3_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_7_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_7_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_7_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_7_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_7_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_7_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_7_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_7_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_7_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_7_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_7_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_7_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_7_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_7_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_7_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_7_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_7_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_7_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_3_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_3_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_3_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_3_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_3_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_3_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_3_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_3_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_3_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_3_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_3_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_3_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_3_norm2_HAS_BIAS = 1,
    parameter stream_blocks_3_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_3_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_3_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_3_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_3_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_3_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_3_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_3_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_3_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_3_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_3_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_3_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_3_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_8_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_8_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_8_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_8_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_8_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_8_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_8_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_8_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_8_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_8_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_8_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_8_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_8_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_8_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_8_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_8_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_8_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_8_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_4_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_4_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_4_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_4_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_4_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_4_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_4_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_4_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_4_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_4_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_4_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_4_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_4_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_4_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_4_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_4_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_4_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_4_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_4_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_4_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_4_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_4_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_4_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_4_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_4_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_4_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_4_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_4_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_4_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_4_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_4_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_4_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_4_norm1_HAS_BIAS = 1,
    parameter stream_blocks_4_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_4_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_4_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_4_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_4_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_4_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_4_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_4_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_4_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_9_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_9_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_9_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_9_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_9_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_9_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_9_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_9_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_9_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_9_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_9_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_9_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_9_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_9_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_9_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_9_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_9_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_9_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_4_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_4_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_4_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_4_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_4_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_4_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_4_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_4_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_4_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_4_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_4_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_4_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_4_norm2_HAS_BIAS = 1,
    parameter stream_blocks_4_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_4_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_4_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_4_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_4_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_4_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_4_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_4_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_4_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_4_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_4_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_4_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_4_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_10_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_10_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_10_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_10_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_10_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_10_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_10_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_10_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_10_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_10_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_10_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_10_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_10_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_10_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_10_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_10_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_10_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_10_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_5_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_5_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_5_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_5_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_5_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_5_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_5_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_5_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_5_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_5_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_5_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_5_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_5_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_5_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_5_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_5_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_5_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_5_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_5_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_5_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_5_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_5_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_5_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_5_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_5_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_5_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_5_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_5_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_5_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_5_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_5_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_5_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_5_norm1_HAS_BIAS = 1,
    parameter stream_blocks_5_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_5_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_5_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_5_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_5_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_5_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_5_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_5_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_5_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_11_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_11_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_11_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_11_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_11_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_11_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_11_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_11_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_11_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_11_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_11_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_11_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_11_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_11_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_11_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_11_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_11_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_11_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_5_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_5_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_5_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_5_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_5_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_5_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_5_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_5_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_5_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_5_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_5_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_5_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_5_norm2_HAS_BIAS = 1,
    parameter stream_blocks_5_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_5_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_5_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_5_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_5_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_5_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_5_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_5_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_5_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_5_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_5_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_5_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_5_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_12_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_12_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_12_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_12_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_12_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_12_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_12_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_12_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_12_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_12_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_12_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_12_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_12_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_12_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_12_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_12_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_12_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_12_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_6_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_6_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_6_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_6_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_6_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_6_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_6_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_6_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_6_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_6_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_6_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_6_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_6_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_6_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_6_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_6_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_6_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_6_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_6_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_6_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_6_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_6_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_6_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_6_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_6_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_6_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_6_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_6_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_6_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_6_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_6_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_6_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_6_norm1_HAS_BIAS = 1,
    parameter stream_blocks_6_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_6_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_6_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_6_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_6_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_6_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_6_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_6_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_6_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_13_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_13_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_13_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_13_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_13_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_13_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_13_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_13_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_13_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_13_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_13_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_13_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_13_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_13_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_13_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_13_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_13_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_13_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_6_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_6_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_6_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_6_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_6_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_6_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_6_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_6_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_6_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_6_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_6_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_6_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_6_norm2_HAS_BIAS = 1,
    parameter stream_blocks_6_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_6_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_6_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_6_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_6_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_6_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_6_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_6_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_6_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_6_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_6_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_6_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_6_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_14_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_14_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_14_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_14_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_14_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_14_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_14_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_14_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_14_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_14_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_14_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_14_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_14_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_14_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_14_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_14_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_14_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_14_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_7_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_7_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_7_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_7_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_7_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_7_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_7_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_7_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_7_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_7_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_7_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_7_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_7_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_7_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_7_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_7_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_7_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_7_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_7_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_7_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_7_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_7_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_7_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_7_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_7_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_7_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_7_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_7_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_7_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_7_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_7_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_7_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_7_norm1_HAS_BIAS = 1,
    parameter stream_blocks_7_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_7_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_7_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_7_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_7_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_7_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_7_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_7_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_7_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_15_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_15_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_15_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_15_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_15_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_15_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_15_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_15_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_15_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_15_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_15_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_15_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_15_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_15_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_15_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_15_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_15_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_15_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_7_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_7_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_7_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_7_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_7_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_7_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_7_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_7_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_7_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_7_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_7_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_7_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_7_norm2_HAS_BIAS = 1,
    parameter stream_blocks_7_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_7_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_7_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_7_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_7_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_7_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_7_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_7_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_7_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_7_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_7_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_7_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_7_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_16_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_16_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_16_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_16_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_16_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_16_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_16_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_16_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_16_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_16_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_16_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_16_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_16_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_16_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_16_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_16_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_16_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_16_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_8_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_8_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_8_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_8_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_8_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_8_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_8_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_8_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_8_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_8_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_8_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_8_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_8_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_8_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_8_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_8_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_8_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_8_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_8_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_8_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_8_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_8_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_8_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_8_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_8_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_8_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_8_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_8_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_8_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_8_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_8_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_8_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_8_norm1_HAS_BIAS = 1,
    parameter stream_blocks_8_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_8_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_8_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_8_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_8_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_8_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_8_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_8_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_8_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_17_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_17_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_17_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_17_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_17_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_17_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_17_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_17_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_17_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_17_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_17_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_17_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_17_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_17_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_17_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_17_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_17_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_17_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_8_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_8_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_8_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_8_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_8_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_8_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_8_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_8_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_8_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_8_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_8_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_8_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_8_norm2_HAS_BIAS = 1,
    parameter stream_blocks_8_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_8_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_8_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_8_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_8_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_8_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_8_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_8_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_8_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_8_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_8_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_8_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_8_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_18_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_18_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_18_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_18_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_18_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_18_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_18_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_18_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_18_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_18_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_18_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_18_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_18_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_18_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_18_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_18_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_18_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_18_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_9_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_9_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_9_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_9_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_9_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_9_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_9_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_9_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_9_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_9_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_9_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_9_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_9_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_9_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_9_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_9_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_9_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_9_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_9_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_9_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_9_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_9_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_9_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_9_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_9_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_9_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_9_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_9_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_9_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_9_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_9_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_9_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_9_norm1_HAS_BIAS = 1,
    parameter stream_blocks_9_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_9_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_9_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_9_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_9_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_9_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_9_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_9_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_9_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_19_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_19_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_19_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_19_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_19_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_19_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_19_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_19_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_19_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_19_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_19_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_19_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_19_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_19_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_19_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_19_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_19_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_19_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_9_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_9_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_9_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_9_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_9_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_9_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_9_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_9_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_9_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_9_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_9_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_9_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_9_norm2_HAS_BIAS = 1,
    parameter stream_blocks_9_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_9_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_9_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_9_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_9_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_9_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_9_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_9_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_9_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_9_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_9_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_9_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_9_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_20_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_20_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_20_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_20_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_20_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_20_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_20_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_20_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_20_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_20_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_20_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_20_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_20_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_20_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_20_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_20_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_20_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_20_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_10_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_10_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_10_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_10_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_10_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_10_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_10_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_10_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_10_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_10_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_10_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_10_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_10_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_10_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_10_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_10_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_10_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_10_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_10_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_10_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_10_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_10_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_10_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_10_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_10_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_10_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_10_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_10_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_10_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_10_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_10_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_10_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_10_norm1_HAS_BIAS = 1,
    parameter stream_blocks_10_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_10_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_10_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_10_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_10_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_10_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_10_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_10_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_10_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_21_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_21_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_21_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_21_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_21_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_21_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_21_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_21_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_21_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_21_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_21_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_21_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_21_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_21_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_21_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_21_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_21_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_21_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_10_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_10_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_10_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_10_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_10_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_10_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_10_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_10_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_10_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_10_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_10_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_10_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_10_norm2_HAS_BIAS = 1,
    parameter stream_blocks_10_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_10_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_10_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_10_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_10_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_10_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_10_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_10_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_10_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_10_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_10_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_10_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_10_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_22_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_22_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_22_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_22_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_22_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_22_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_22_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_22_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_22_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_22_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_22_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_22_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_22_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_22_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_22_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_22_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_22_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_22_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_linear1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_11_linear1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_11_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_linear1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_linear1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_linear1_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_11_linear1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_11_linear1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_linear1_WEIGHT_TENSOR_SIZE_DIM_1 = 768,
    parameter stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_11_linear1_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_11_linear1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_11_linear1_BIAS_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_linear1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_linear1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_11_linear1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_11_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_11_linear1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_linear1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_act_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_11_act_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_11_act_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_11_act_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_act_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_act_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_act_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_11_act_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_11_act_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_11_act_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_act_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_act_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_linear2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_11_linear2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_11_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_11_linear2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_linear2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_linear2_WEIGHT_PRECISION_0 = 4,
    parameter stream_blocks_11_linear2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_11_linear2_WEIGHT_TENSOR_SIZE_DIM_0 = 768,
    parameter stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_linear2_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_11_linear2_BIAS_PRECISION_0 = 4,
    parameter stream_blocks_11_linear2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_11_linear2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_linear2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_linear2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_11_linear2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_11_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_linear2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_linear2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_norm1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_11_norm1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_11_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_norm1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_norm1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_norm1_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_11_norm1_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_11_norm1_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_norm1_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_norm1_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_11_norm1_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_11_norm1_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_norm1_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_norm1_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_11_norm1_HAS_BIAS = 1,
    parameter stream_blocks_11_norm1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_11_norm1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_11_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_norm1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_norm1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_add_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_11_add_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_11_add_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_add_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_add_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_add_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_add_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_11_add_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_11_add_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_add_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_add_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_add_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_add_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_11_add_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_11_add_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_add_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_add_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_add_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_23_DATA_IN_0_PRECISION_0 = 6,
    parameter fork2_23_DATA_IN_0_PRECISION_1 = 4,
    parameter fork2_23_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_23_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_23_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_23_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_23_DATA_OUT_0_PRECISION_0 = 6,
    parameter fork2_23_DATA_OUT_0_PRECISION_1 = 4,
    parameter fork2_23_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_23_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter fork2_23_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_23_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter fork2_23_DATA_OUT_1_PRECISION_0 = 6,
    parameter fork2_23_DATA_OUT_1_PRECISION_1 = 4,
    parameter fork2_23_DATA_OUT_1_TENSOR_SIZE_DIM_0 = 192,
    parameter fork2_23_DATA_OUT_1_PARALLELISM_DIM_0 = 4,
    parameter fork2_23_DATA_OUT_1_TENSOR_SIZE_DIM_1 = 196,
    parameter fork2_23_DATA_OUT_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_attention_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_attention_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_11_attention_QUERY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_QUERY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_attention_KEY_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_KEY_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_11_attention_KEY_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_KEY_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_KEY_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_KEY_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_11_attention_VALUE_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_VALUE_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1 = 192,
    parameter stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_1 = 4,
    parameter stream_blocks_11_attention_PROJ_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_PROJ_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_attention_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_11_attention_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_11_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_attention_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_attention_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_norm2_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_11_norm2_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_11_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_norm2_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_norm2_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_norm2_WEIGHT_PRECISION_0 = 6,
    parameter stream_blocks_11_norm2_WEIGHT_PRECISION_1 = 4,
    parameter stream_blocks_11_norm2_WEIGHT_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_norm2_WEIGHT_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_norm2_BIAS_PRECISION_0 = 6,
    parameter stream_blocks_11_norm2_BIAS_PRECISION_1 = 4,
    parameter stream_blocks_11_norm2_BIAS_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_norm2_BIAS_TENSOR_SIZE_DIM_1 = 1,
    parameter stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_norm2_ELEMENTWISE_AFFINE = 1,
    parameter stream_blocks_11_norm2_HAS_BIAS = 1,
    parameter stream_blocks_11_norm2_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_11_norm2_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_11_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_norm2_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_norm2_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_add_1_DATA_IN_0_PRECISION_0 = 6,
    parameter stream_blocks_11_add_1_DATA_IN_0_PRECISION_1 = 4,
    parameter stream_blocks_11_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_add_1_DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_add_1_DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_add_1_DATA_IN_1_PRECISION_0 = 6,
    parameter stream_blocks_11_add_1_DATA_IN_1_PRECISION_1 = 4,
    parameter stream_blocks_11_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_add_1_DATA_IN_1_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_add_1_DATA_IN_1_PARALLELISM_DIM_1 = 1,
    parameter stream_blocks_11_add_1_DATA_OUT_0_PRECISION_0 = 6,
    parameter stream_blocks_11_add_1_DATA_OUT_0_PRECISION_1 = 4,
    parameter stream_blocks_11_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter stream_blocks_11_add_1_DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter stream_blocks_11_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter stream_blocks_11_add_1_DATA_OUT_0_PARALLELISM_DIM_1 = 1,
    parameter DATA_IN_0_PRECISION_0 = 6,
    parameter DATA_IN_0_PRECISION_1 = 4,
    parameter DATA_IN_0_TENSOR_SIZE_DIM_0 = 192,
    parameter DATA_IN_0_PARALLELISM_DIM_0 = 4,
    parameter DATA_IN_0_TENSOR_SIZE_DIM_1 = 196,
    parameter DATA_IN_0_PARALLELISM_DIM_1 = 1,
    parameter DATA_OUT_0_PRECISION_0 = 6,
    parameter DATA_OUT_0_PRECISION_1 = 4,
    parameter DATA_OUT_0_TENSOR_SIZE_DIM_0 = 192,
    parameter DATA_OUT_0_PARALLELISM_DIM_0 = 4,
    parameter DATA_OUT_0_TENSOR_SIZE_DIM_1 = 196,
    parameter DATA_OUT_0_PARALLELISM_DIM_1 = 1
) (
    input clk,
    input rst,

    input  [DATA_IN_0_PRECISION_0-1:0] mdata_in_0 [DATA_IN_0_PARALLELISM_DIM_0*DATA_IN_0_PARALLELISM_DIM_1-1:0],
    input  [DATA_IN_0_PRECISION_1-1:0] edata_in_0,
    input  data_in_0_valid,
    output data_in_0_ready,
    output  [DATA_OUT_0_PRECISION_0-1:0] mdata_out_0 [DATA_OUT_0_PARALLELISM_DIM_0*DATA_OUT_0_PARALLELISM_DIM_1-1:0],
    output  [DATA_OUT_0_PRECISION_1-1:0] edata_out_0,
    output  data_out_0_valid,
    input data_out_0_ready
);

// --------------------------
//   fork2 signals
// --------------------------
logic [fork2_DATA_IN_0_PRECISION_0-1:0]  fork2_mdata_in_0        [fork2_DATA_IN_0_PARALLELISM_DIM_0*fork2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_DATA_IN_0_PRECISION_1-1:0]  fork2_edata_in_0;
logic                             fork2_data_in_0_valid;
logic                             fork2_data_in_0_ready;
logic [fork2_DATA_OUT_0_PRECISION_0-1:0]  fork2_mdata_out_0        [fork2_DATA_OUT_0_PARALLELISM_DIM_0*fork2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_DATA_OUT_0_PRECISION_1-1:0]  fork2_edata_out_0;
logic                             fork2_data_out_0_valid;
logic                             fork2_data_out_0_ready;
logic [fork2_DATA_OUT_1_PRECISION_0-1:0]  fork2_mdata_out_1        [fork2_DATA_OUT_1_PARALLELISM_DIM_0*fork2_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_DATA_OUT_1_PRECISION_1-1:0]  fork2_edata_out_1;
logic                             fork2_data_out_1_valid;
logic                             fork2_data_out_1_ready;
// --------------------------
//   stream_blocks_0_linear1 signals
// --------------------------
logic [stream_blocks_0_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_0_linear1_mdata_in_0        [stream_blocks_0_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_0_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_0_linear1_edata_in_0;
logic                             stream_blocks_0_linear1_data_in_0_valid;
logic                             stream_blocks_0_linear1_data_in_0_ready;
logic [stream_blocks_0_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_0_linear1_mweight        [stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_0_linear1_eweight;
logic                             stream_blocks_0_linear1_weight_valid;
logic                             stream_blocks_0_linear1_weight_ready;
logic [stream_blocks_0_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_0_linear1_mbias        [stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_0_linear1_ebias;
logic                             stream_blocks_0_linear1_bias_valid;
logic                             stream_blocks_0_linear1_bias_ready;
logic [stream_blocks_0_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_0_linear1_mdata_out_0        [stream_blocks_0_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_0_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_0_linear1_edata_out_0;
logic                             stream_blocks_0_linear1_data_out_0_valid;
logic                             stream_blocks_0_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_0_act signals
// --------------------------
logic [stream_blocks_0_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_0_act_mdata_in_0        [stream_blocks_0_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_0_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_0_act_edata_in_0;
logic                             stream_blocks_0_act_data_in_0_valid;
logic                             stream_blocks_0_act_data_in_0_ready;
logic [stream_blocks_0_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_0_act_mdata_out_0        [stream_blocks_0_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_0_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_0_act_edata_out_0;
logic                             stream_blocks_0_act_data_out_0_valid;
logic                             stream_blocks_0_act_data_out_0_ready;
// --------------------------
//   stream_blocks_0_linear2 signals
// --------------------------
logic [stream_blocks_0_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_0_linear2_mdata_in_0        [stream_blocks_0_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_0_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_0_linear2_edata_in_0;
logic                             stream_blocks_0_linear2_data_in_0_valid;
logic                             stream_blocks_0_linear2_data_in_0_ready;
logic [stream_blocks_0_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_0_linear2_mweight        [stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_0_linear2_eweight;
logic                             stream_blocks_0_linear2_weight_valid;
logic                             stream_blocks_0_linear2_weight_ready;
logic [stream_blocks_0_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_0_linear2_mbias        [stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_0_linear2_ebias;
logic                             stream_blocks_0_linear2_bias_valid;
logic                             stream_blocks_0_linear2_bias_ready;
logic [stream_blocks_0_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_0_linear2_mdata_out_0        [stream_blocks_0_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_0_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_0_linear2_edata_out_0;
logic                             stream_blocks_0_linear2_data_out_0_valid;
logic                             stream_blocks_0_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_0_norm1 signals
// --------------------------
logic [stream_blocks_0_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_0_norm1_mdata_in_0        [stream_blocks_0_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_0_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_0_norm1_edata_in_0;
logic                             stream_blocks_0_norm1_data_in_0_valid;
logic                             stream_blocks_0_norm1_data_in_0_ready;
logic [stream_blocks_0_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_0_norm1_mweight        [stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_0_norm1_eweight;
logic                             stream_blocks_0_norm1_weight_valid;
logic                             stream_blocks_0_norm1_weight_ready;
logic [stream_blocks_0_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_0_norm1_mbias        [stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_0_norm1_ebias;
logic                             stream_blocks_0_norm1_bias_valid;
logic                             stream_blocks_0_norm1_bias_ready;
logic [stream_blocks_0_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_0_norm1_mdata_out_0        [stream_blocks_0_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_0_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_0_norm1_edata_out_0;
logic                             stream_blocks_0_norm1_data_out_0_valid;
logic                             stream_blocks_0_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_0_add signals
// --------------------------
logic [stream_blocks_0_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_0_add_mdata_in_0        [stream_blocks_0_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_0_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_0_add_edata_in_0;
logic                             stream_blocks_0_add_data_in_0_valid;
logic                             stream_blocks_0_add_data_in_0_ready;
logic [stream_blocks_0_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_0_add_mdata_in_1        [stream_blocks_0_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_0_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_0_add_edata_in_1;
logic                             stream_blocks_0_add_data_in_1_valid;
logic                             stream_blocks_0_add_data_in_1_ready;
logic [stream_blocks_0_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_0_add_mdata_out_0        [stream_blocks_0_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_0_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_0_add_edata_out_0;
logic                             stream_blocks_0_add_data_out_0_valid;
logic                             stream_blocks_0_add_data_out_0_ready;
// --------------------------
//   fork2_1 signals
// --------------------------
logic [fork2_1_DATA_IN_0_PRECISION_0-1:0]  fork2_1_mdata_in_0        [fork2_1_DATA_IN_0_PARALLELISM_DIM_0*fork2_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_1_DATA_IN_0_PRECISION_1-1:0]  fork2_1_edata_in_0;
logic                             fork2_1_data_in_0_valid;
logic                             fork2_1_data_in_0_ready;
logic [fork2_1_DATA_OUT_0_PRECISION_0-1:0]  fork2_1_mdata_out_0        [fork2_1_DATA_OUT_0_PARALLELISM_DIM_0*fork2_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_1_DATA_OUT_0_PRECISION_1-1:0]  fork2_1_edata_out_0;
logic                             fork2_1_data_out_0_valid;
logic                             fork2_1_data_out_0_ready;
logic [fork2_1_DATA_OUT_1_PRECISION_0-1:0]  fork2_1_mdata_out_1        [fork2_1_DATA_OUT_1_PARALLELISM_DIM_0*fork2_1_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_1_DATA_OUT_1_PRECISION_1-1:0]  fork2_1_edata_out_1;
logic                             fork2_1_data_out_1_valid;
logic                             fork2_1_data_out_1_ready;
// --------------------------
//   stream_blocks_0_attention signals
// --------------------------
logic [stream_blocks_0_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_0_attention_mdata_in_0        [stream_blocks_0_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_0_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_0_attention_edata_in_0;
logic                             stream_blocks_0_attention_data_in_0_valid;
logic                             stream_blocks_0_attention_data_in_0_ready;
logic [stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_0_attention_mquery_weight        [stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_0_attention_equery_weight;
logic                             stream_blocks_0_attention_query_weight_valid;
logic                             stream_blocks_0_attention_query_weight_ready;
logic [stream_blocks_0_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_0_attention_mquery_bias        [stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_0_attention_equery_bias;
logic                             stream_blocks_0_attention_query_bias_valid;
logic                             stream_blocks_0_attention_query_bias_ready;
logic [stream_blocks_0_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_0_attention_mkey_weight        [stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_0_attention_ekey_weight;
logic                             stream_blocks_0_attention_key_weight_valid;
logic                             stream_blocks_0_attention_key_weight_ready;
logic [stream_blocks_0_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_0_attention_mkey_bias        [stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_0_attention_ekey_bias;
logic                             stream_blocks_0_attention_key_bias_valid;
logic                             stream_blocks_0_attention_key_bias_ready;
logic [stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_0_attention_mvalue_weight        [stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_0_attention_evalue_weight;
logic                             stream_blocks_0_attention_value_weight_valid;
logic                             stream_blocks_0_attention_value_weight_ready;
logic [stream_blocks_0_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_0_attention_mvalue_bias        [stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_0_attention_evalue_bias;
logic                             stream_blocks_0_attention_value_bias_valid;
logic                             stream_blocks_0_attention_value_bias_ready;
logic [stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_0_attention_mproj_weight        [stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_0_attention_eproj_weight;
logic                             stream_blocks_0_attention_proj_weight_valid;
logic                             stream_blocks_0_attention_proj_weight_ready;
logic [stream_blocks_0_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_0_attention_mproj_bias        [stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_0_attention_eproj_bias;
logic                             stream_blocks_0_attention_proj_bias_valid;
logic                             stream_blocks_0_attention_proj_bias_ready;
logic [stream_blocks_0_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_0_attention_mdata_out_0        [stream_blocks_0_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_0_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_0_attention_edata_out_0;
logic                             stream_blocks_0_attention_data_out_0_valid;
logic                             stream_blocks_0_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_0_norm2 signals
// --------------------------
logic [stream_blocks_0_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_0_norm2_mdata_in_0        [stream_blocks_0_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_0_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_0_norm2_edata_in_0;
logic                             stream_blocks_0_norm2_data_in_0_valid;
logic                             stream_blocks_0_norm2_data_in_0_ready;
logic [stream_blocks_0_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_0_norm2_mweight        [stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_0_norm2_eweight;
logic                             stream_blocks_0_norm2_weight_valid;
logic                             stream_blocks_0_norm2_weight_ready;
logic [stream_blocks_0_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_0_norm2_mbias        [stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_0_norm2_ebias;
logic                             stream_blocks_0_norm2_bias_valid;
logic                             stream_blocks_0_norm2_bias_ready;
logic [stream_blocks_0_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_0_norm2_mdata_out_0        [stream_blocks_0_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_0_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_0_norm2_edata_out_0;
logic                             stream_blocks_0_norm2_data_out_0_valid;
logic                             stream_blocks_0_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_0_add_1 signals
// --------------------------
logic [stream_blocks_0_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_0_add_1_mdata_in_0        [stream_blocks_0_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_0_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_0_add_1_edata_in_0;
logic                             stream_blocks_0_add_1_data_in_0_valid;
logic                             stream_blocks_0_add_1_data_in_0_ready;
logic [stream_blocks_0_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_0_add_1_mdata_in_1        [stream_blocks_0_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_0_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_0_add_1_edata_in_1;
logic                             stream_blocks_0_add_1_data_in_1_valid;
logic                             stream_blocks_0_add_1_data_in_1_ready;
logic [stream_blocks_0_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_0_add_1_mdata_out_0        [stream_blocks_0_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_0_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_0_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_0_add_1_edata_out_0;
logic                             stream_blocks_0_add_1_data_out_0_valid;
logic                             stream_blocks_0_add_1_data_out_0_ready;
// --------------------------
//   fork2_2 signals
// --------------------------
logic [fork2_2_DATA_IN_0_PRECISION_0-1:0]  fork2_2_mdata_in_0        [fork2_2_DATA_IN_0_PARALLELISM_DIM_0*fork2_2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_2_DATA_IN_0_PRECISION_1-1:0]  fork2_2_edata_in_0;
logic                             fork2_2_data_in_0_valid;
logic                             fork2_2_data_in_0_ready;
logic [fork2_2_DATA_OUT_0_PRECISION_0-1:0]  fork2_2_mdata_out_0        [fork2_2_DATA_OUT_0_PARALLELISM_DIM_0*fork2_2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_2_DATA_OUT_0_PRECISION_1-1:0]  fork2_2_edata_out_0;
logic                             fork2_2_data_out_0_valid;
logic                             fork2_2_data_out_0_ready;
logic [fork2_2_DATA_OUT_1_PRECISION_0-1:0]  fork2_2_mdata_out_1        [fork2_2_DATA_OUT_1_PARALLELISM_DIM_0*fork2_2_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_2_DATA_OUT_1_PRECISION_1-1:0]  fork2_2_edata_out_1;
logic                             fork2_2_data_out_1_valid;
logic                             fork2_2_data_out_1_ready;
// --------------------------
//   stream_blocks_1_linear1 signals
// --------------------------
logic [stream_blocks_1_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_1_linear1_mdata_in_0        [stream_blocks_1_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_1_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_1_linear1_edata_in_0;
logic                             stream_blocks_1_linear1_data_in_0_valid;
logic                             stream_blocks_1_linear1_data_in_0_ready;
logic [stream_blocks_1_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_1_linear1_mweight        [stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_1_linear1_eweight;
logic                             stream_blocks_1_linear1_weight_valid;
logic                             stream_blocks_1_linear1_weight_ready;
logic [stream_blocks_1_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_1_linear1_mbias        [stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_1_linear1_ebias;
logic                             stream_blocks_1_linear1_bias_valid;
logic                             stream_blocks_1_linear1_bias_ready;
logic [stream_blocks_1_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_1_linear1_mdata_out_0        [stream_blocks_1_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_1_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_1_linear1_edata_out_0;
logic                             stream_blocks_1_linear1_data_out_0_valid;
logic                             stream_blocks_1_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_1_act signals
// --------------------------
logic [stream_blocks_1_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_1_act_mdata_in_0        [stream_blocks_1_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_1_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_1_act_edata_in_0;
logic                             stream_blocks_1_act_data_in_0_valid;
logic                             stream_blocks_1_act_data_in_0_ready;
logic [stream_blocks_1_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_1_act_mdata_out_0        [stream_blocks_1_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_1_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_1_act_edata_out_0;
logic                             stream_blocks_1_act_data_out_0_valid;
logic                             stream_blocks_1_act_data_out_0_ready;
// --------------------------
//   stream_blocks_1_linear2 signals
// --------------------------
logic [stream_blocks_1_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_1_linear2_mdata_in_0        [stream_blocks_1_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_1_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_1_linear2_edata_in_0;
logic                             stream_blocks_1_linear2_data_in_0_valid;
logic                             stream_blocks_1_linear2_data_in_0_ready;
logic [stream_blocks_1_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_1_linear2_mweight        [stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_1_linear2_eweight;
logic                             stream_blocks_1_linear2_weight_valid;
logic                             stream_blocks_1_linear2_weight_ready;
logic [stream_blocks_1_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_1_linear2_mbias        [stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_1_linear2_ebias;
logic                             stream_blocks_1_linear2_bias_valid;
logic                             stream_blocks_1_linear2_bias_ready;
logic [stream_blocks_1_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_1_linear2_mdata_out_0        [stream_blocks_1_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_1_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_1_linear2_edata_out_0;
logic                             stream_blocks_1_linear2_data_out_0_valid;
logic                             stream_blocks_1_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_1_norm1 signals
// --------------------------
logic [stream_blocks_1_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_1_norm1_mdata_in_0        [stream_blocks_1_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_1_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_1_norm1_edata_in_0;
logic                             stream_blocks_1_norm1_data_in_0_valid;
logic                             stream_blocks_1_norm1_data_in_0_ready;
logic [stream_blocks_1_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_1_norm1_mweight        [stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_1_norm1_eweight;
logic                             stream_blocks_1_norm1_weight_valid;
logic                             stream_blocks_1_norm1_weight_ready;
logic [stream_blocks_1_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_1_norm1_mbias        [stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_1_norm1_ebias;
logic                             stream_blocks_1_norm1_bias_valid;
logic                             stream_blocks_1_norm1_bias_ready;
logic [stream_blocks_1_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_1_norm1_mdata_out_0        [stream_blocks_1_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_1_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_1_norm1_edata_out_0;
logic                             stream_blocks_1_norm1_data_out_0_valid;
logic                             stream_blocks_1_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_1_add signals
// --------------------------
logic [stream_blocks_1_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_1_add_mdata_in_0        [stream_blocks_1_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_1_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_1_add_edata_in_0;
logic                             stream_blocks_1_add_data_in_0_valid;
logic                             stream_blocks_1_add_data_in_0_ready;
logic [stream_blocks_1_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_1_add_mdata_in_1        [stream_blocks_1_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_1_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_1_add_edata_in_1;
logic                             stream_blocks_1_add_data_in_1_valid;
logic                             stream_blocks_1_add_data_in_1_ready;
logic [stream_blocks_1_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_1_add_mdata_out_0        [stream_blocks_1_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_1_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_1_add_edata_out_0;
logic                             stream_blocks_1_add_data_out_0_valid;
logic                             stream_blocks_1_add_data_out_0_ready;
// --------------------------
//   fork2_3 signals
// --------------------------
logic [fork2_3_DATA_IN_0_PRECISION_0-1:0]  fork2_3_mdata_in_0        [fork2_3_DATA_IN_0_PARALLELISM_DIM_0*fork2_3_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_3_DATA_IN_0_PRECISION_1-1:0]  fork2_3_edata_in_0;
logic                             fork2_3_data_in_0_valid;
logic                             fork2_3_data_in_0_ready;
logic [fork2_3_DATA_OUT_0_PRECISION_0-1:0]  fork2_3_mdata_out_0        [fork2_3_DATA_OUT_0_PARALLELISM_DIM_0*fork2_3_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_3_DATA_OUT_0_PRECISION_1-1:0]  fork2_3_edata_out_0;
logic                             fork2_3_data_out_0_valid;
logic                             fork2_3_data_out_0_ready;
logic [fork2_3_DATA_OUT_1_PRECISION_0-1:0]  fork2_3_mdata_out_1        [fork2_3_DATA_OUT_1_PARALLELISM_DIM_0*fork2_3_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_3_DATA_OUT_1_PRECISION_1-1:0]  fork2_3_edata_out_1;
logic                             fork2_3_data_out_1_valid;
logic                             fork2_3_data_out_1_ready;
// --------------------------
//   stream_blocks_1_attention signals
// --------------------------
logic [stream_blocks_1_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_1_attention_mdata_in_0        [stream_blocks_1_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_1_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_1_attention_edata_in_0;
logic                             stream_blocks_1_attention_data_in_0_valid;
logic                             stream_blocks_1_attention_data_in_0_ready;
logic [stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_1_attention_mquery_weight        [stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_1_attention_equery_weight;
logic                             stream_blocks_1_attention_query_weight_valid;
logic                             stream_blocks_1_attention_query_weight_ready;
logic [stream_blocks_1_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_1_attention_mquery_bias        [stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_1_attention_equery_bias;
logic                             stream_blocks_1_attention_query_bias_valid;
logic                             stream_blocks_1_attention_query_bias_ready;
logic [stream_blocks_1_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_1_attention_mkey_weight        [stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_1_attention_ekey_weight;
logic                             stream_blocks_1_attention_key_weight_valid;
logic                             stream_blocks_1_attention_key_weight_ready;
logic [stream_blocks_1_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_1_attention_mkey_bias        [stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_1_attention_ekey_bias;
logic                             stream_blocks_1_attention_key_bias_valid;
logic                             stream_blocks_1_attention_key_bias_ready;
logic [stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_1_attention_mvalue_weight        [stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_1_attention_evalue_weight;
logic                             stream_blocks_1_attention_value_weight_valid;
logic                             stream_blocks_1_attention_value_weight_ready;
logic [stream_blocks_1_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_1_attention_mvalue_bias        [stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_1_attention_evalue_bias;
logic                             stream_blocks_1_attention_value_bias_valid;
logic                             stream_blocks_1_attention_value_bias_ready;
logic [stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_1_attention_mproj_weight        [stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_1_attention_eproj_weight;
logic                             stream_blocks_1_attention_proj_weight_valid;
logic                             stream_blocks_1_attention_proj_weight_ready;
logic [stream_blocks_1_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_1_attention_mproj_bias        [stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_1_attention_eproj_bias;
logic                             stream_blocks_1_attention_proj_bias_valid;
logic                             stream_blocks_1_attention_proj_bias_ready;
logic [stream_blocks_1_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_1_attention_mdata_out_0        [stream_blocks_1_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_1_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_1_attention_edata_out_0;
logic                             stream_blocks_1_attention_data_out_0_valid;
logic                             stream_blocks_1_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_1_norm2 signals
// --------------------------
logic [stream_blocks_1_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_1_norm2_mdata_in_0        [stream_blocks_1_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_1_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_1_norm2_edata_in_0;
logic                             stream_blocks_1_norm2_data_in_0_valid;
logic                             stream_blocks_1_norm2_data_in_0_ready;
logic [stream_blocks_1_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_1_norm2_mweight        [stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_1_norm2_eweight;
logic                             stream_blocks_1_norm2_weight_valid;
logic                             stream_blocks_1_norm2_weight_ready;
logic [stream_blocks_1_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_1_norm2_mbias        [stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_1_norm2_ebias;
logic                             stream_blocks_1_norm2_bias_valid;
logic                             stream_blocks_1_norm2_bias_ready;
logic [stream_blocks_1_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_1_norm2_mdata_out_0        [stream_blocks_1_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_1_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_1_norm2_edata_out_0;
logic                             stream_blocks_1_norm2_data_out_0_valid;
logic                             stream_blocks_1_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_1_add_1 signals
// --------------------------
logic [stream_blocks_1_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_1_add_1_mdata_in_0        [stream_blocks_1_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_1_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_1_add_1_edata_in_0;
logic                             stream_blocks_1_add_1_data_in_0_valid;
logic                             stream_blocks_1_add_1_data_in_0_ready;
logic [stream_blocks_1_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_1_add_1_mdata_in_1        [stream_blocks_1_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_1_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_1_add_1_edata_in_1;
logic                             stream_blocks_1_add_1_data_in_1_valid;
logic                             stream_blocks_1_add_1_data_in_1_ready;
logic [stream_blocks_1_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_1_add_1_mdata_out_0        [stream_blocks_1_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_1_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_1_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_1_add_1_edata_out_0;
logic                             stream_blocks_1_add_1_data_out_0_valid;
logic                             stream_blocks_1_add_1_data_out_0_ready;
// --------------------------
//   fork2_4 signals
// --------------------------
logic [fork2_4_DATA_IN_0_PRECISION_0-1:0]  fork2_4_mdata_in_0        [fork2_4_DATA_IN_0_PARALLELISM_DIM_0*fork2_4_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_4_DATA_IN_0_PRECISION_1-1:0]  fork2_4_edata_in_0;
logic                             fork2_4_data_in_0_valid;
logic                             fork2_4_data_in_0_ready;
logic [fork2_4_DATA_OUT_0_PRECISION_0-1:0]  fork2_4_mdata_out_0        [fork2_4_DATA_OUT_0_PARALLELISM_DIM_0*fork2_4_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_4_DATA_OUT_0_PRECISION_1-1:0]  fork2_4_edata_out_0;
logic                             fork2_4_data_out_0_valid;
logic                             fork2_4_data_out_0_ready;
logic [fork2_4_DATA_OUT_1_PRECISION_0-1:0]  fork2_4_mdata_out_1        [fork2_4_DATA_OUT_1_PARALLELISM_DIM_0*fork2_4_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_4_DATA_OUT_1_PRECISION_1-1:0]  fork2_4_edata_out_1;
logic                             fork2_4_data_out_1_valid;
logic                             fork2_4_data_out_1_ready;
// --------------------------
//   stream_blocks_2_linear1 signals
// --------------------------
logic [stream_blocks_2_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_2_linear1_mdata_in_0        [stream_blocks_2_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_2_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_2_linear1_edata_in_0;
logic                             stream_blocks_2_linear1_data_in_0_valid;
logic                             stream_blocks_2_linear1_data_in_0_ready;
logic [stream_blocks_2_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_2_linear1_mweight        [stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_2_linear1_eweight;
logic                             stream_blocks_2_linear1_weight_valid;
logic                             stream_blocks_2_linear1_weight_ready;
logic [stream_blocks_2_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_2_linear1_mbias        [stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_2_linear1_ebias;
logic                             stream_blocks_2_linear1_bias_valid;
logic                             stream_blocks_2_linear1_bias_ready;
logic [stream_blocks_2_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_2_linear1_mdata_out_0        [stream_blocks_2_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_2_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_2_linear1_edata_out_0;
logic                             stream_blocks_2_linear1_data_out_0_valid;
logic                             stream_blocks_2_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_2_act signals
// --------------------------
logic [stream_blocks_2_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_2_act_mdata_in_0        [stream_blocks_2_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_2_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_2_act_edata_in_0;
logic                             stream_blocks_2_act_data_in_0_valid;
logic                             stream_blocks_2_act_data_in_0_ready;
logic [stream_blocks_2_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_2_act_mdata_out_0        [stream_blocks_2_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_2_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_2_act_edata_out_0;
logic                             stream_blocks_2_act_data_out_0_valid;
logic                             stream_blocks_2_act_data_out_0_ready;
// --------------------------
//   stream_blocks_2_linear2 signals
// --------------------------
logic [stream_blocks_2_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_2_linear2_mdata_in_0        [stream_blocks_2_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_2_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_2_linear2_edata_in_0;
logic                             stream_blocks_2_linear2_data_in_0_valid;
logic                             stream_blocks_2_linear2_data_in_0_ready;
logic [stream_blocks_2_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_2_linear2_mweight        [stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_2_linear2_eweight;
logic                             stream_blocks_2_linear2_weight_valid;
logic                             stream_blocks_2_linear2_weight_ready;
logic [stream_blocks_2_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_2_linear2_mbias        [stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_2_linear2_ebias;
logic                             stream_blocks_2_linear2_bias_valid;
logic                             stream_blocks_2_linear2_bias_ready;
logic [stream_blocks_2_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_2_linear2_mdata_out_0        [stream_blocks_2_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_2_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_2_linear2_edata_out_0;
logic                             stream_blocks_2_linear2_data_out_0_valid;
logic                             stream_blocks_2_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_2_norm1 signals
// --------------------------
logic [stream_blocks_2_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_2_norm1_mdata_in_0        [stream_blocks_2_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_2_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_2_norm1_edata_in_0;
logic                             stream_blocks_2_norm1_data_in_0_valid;
logic                             stream_blocks_2_norm1_data_in_0_ready;
logic [stream_blocks_2_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_2_norm1_mweight        [stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_2_norm1_eweight;
logic                             stream_blocks_2_norm1_weight_valid;
logic                             stream_blocks_2_norm1_weight_ready;
logic [stream_blocks_2_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_2_norm1_mbias        [stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_2_norm1_ebias;
logic                             stream_blocks_2_norm1_bias_valid;
logic                             stream_blocks_2_norm1_bias_ready;
logic [stream_blocks_2_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_2_norm1_mdata_out_0        [stream_blocks_2_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_2_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_2_norm1_edata_out_0;
logic                             stream_blocks_2_norm1_data_out_0_valid;
logic                             stream_blocks_2_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_2_add signals
// --------------------------
logic [stream_blocks_2_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_2_add_mdata_in_0        [stream_blocks_2_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_2_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_2_add_edata_in_0;
logic                             stream_blocks_2_add_data_in_0_valid;
logic                             stream_blocks_2_add_data_in_0_ready;
logic [stream_blocks_2_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_2_add_mdata_in_1        [stream_blocks_2_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_2_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_2_add_edata_in_1;
logic                             stream_blocks_2_add_data_in_1_valid;
logic                             stream_blocks_2_add_data_in_1_ready;
logic [stream_blocks_2_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_2_add_mdata_out_0        [stream_blocks_2_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_2_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_2_add_edata_out_0;
logic                             stream_blocks_2_add_data_out_0_valid;
logic                             stream_blocks_2_add_data_out_0_ready;
// --------------------------
//   fork2_5 signals
// --------------------------
logic [fork2_5_DATA_IN_0_PRECISION_0-1:0]  fork2_5_mdata_in_0        [fork2_5_DATA_IN_0_PARALLELISM_DIM_0*fork2_5_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_5_DATA_IN_0_PRECISION_1-1:0]  fork2_5_edata_in_0;
logic                             fork2_5_data_in_0_valid;
logic                             fork2_5_data_in_0_ready;
logic [fork2_5_DATA_OUT_0_PRECISION_0-1:0]  fork2_5_mdata_out_0        [fork2_5_DATA_OUT_0_PARALLELISM_DIM_0*fork2_5_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_5_DATA_OUT_0_PRECISION_1-1:0]  fork2_5_edata_out_0;
logic                             fork2_5_data_out_0_valid;
logic                             fork2_5_data_out_0_ready;
logic [fork2_5_DATA_OUT_1_PRECISION_0-1:0]  fork2_5_mdata_out_1        [fork2_5_DATA_OUT_1_PARALLELISM_DIM_0*fork2_5_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_5_DATA_OUT_1_PRECISION_1-1:0]  fork2_5_edata_out_1;
logic                             fork2_5_data_out_1_valid;
logic                             fork2_5_data_out_1_ready;
// --------------------------
//   stream_blocks_2_attention signals
// --------------------------
logic [stream_blocks_2_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_2_attention_mdata_in_0        [stream_blocks_2_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_2_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_2_attention_edata_in_0;
logic                             stream_blocks_2_attention_data_in_0_valid;
logic                             stream_blocks_2_attention_data_in_0_ready;
logic [stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_2_attention_mquery_weight        [stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_2_attention_equery_weight;
logic                             stream_blocks_2_attention_query_weight_valid;
logic                             stream_blocks_2_attention_query_weight_ready;
logic [stream_blocks_2_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_2_attention_mquery_bias        [stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_2_attention_equery_bias;
logic                             stream_blocks_2_attention_query_bias_valid;
logic                             stream_blocks_2_attention_query_bias_ready;
logic [stream_blocks_2_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_2_attention_mkey_weight        [stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_2_attention_ekey_weight;
logic                             stream_blocks_2_attention_key_weight_valid;
logic                             stream_blocks_2_attention_key_weight_ready;
logic [stream_blocks_2_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_2_attention_mkey_bias        [stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_2_attention_ekey_bias;
logic                             stream_blocks_2_attention_key_bias_valid;
logic                             stream_blocks_2_attention_key_bias_ready;
logic [stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_2_attention_mvalue_weight        [stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_2_attention_evalue_weight;
logic                             stream_blocks_2_attention_value_weight_valid;
logic                             stream_blocks_2_attention_value_weight_ready;
logic [stream_blocks_2_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_2_attention_mvalue_bias        [stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_2_attention_evalue_bias;
logic                             stream_blocks_2_attention_value_bias_valid;
logic                             stream_blocks_2_attention_value_bias_ready;
logic [stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_2_attention_mproj_weight        [stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_2_attention_eproj_weight;
logic                             stream_blocks_2_attention_proj_weight_valid;
logic                             stream_blocks_2_attention_proj_weight_ready;
logic [stream_blocks_2_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_2_attention_mproj_bias        [stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_2_attention_eproj_bias;
logic                             stream_blocks_2_attention_proj_bias_valid;
logic                             stream_blocks_2_attention_proj_bias_ready;
logic [stream_blocks_2_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_2_attention_mdata_out_0        [stream_blocks_2_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_2_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_2_attention_edata_out_0;
logic                             stream_blocks_2_attention_data_out_0_valid;
logic                             stream_blocks_2_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_2_norm2 signals
// --------------------------
logic [stream_blocks_2_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_2_norm2_mdata_in_0        [stream_blocks_2_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_2_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_2_norm2_edata_in_0;
logic                             stream_blocks_2_norm2_data_in_0_valid;
logic                             stream_blocks_2_norm2_data_in_0_ready;
logic [stream_blocks_2_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_2_norm2_mweight        [stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_2_norm2_eweight;
logic                             stream_blocks_2_norm2_weight_valid;
logic                             stream_blocks_2_norm2_weight_ready;
logic [stream_blocks_2_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_2_norm2_mbias        [stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_2_norm2_ebias;
logic                             stream_blocks_2_norm2_bias_valid;
logic                             stream_blocks_2_norm2_bias_ready;
logic [stream_blocks_2_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_2_norm2_mdata_out_0        [stream_blocks_2_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_2_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_2_norm2_edata_out_0;
logic                             stream_blocks_2_norm2_data_out_0_valid;
logic                             stream_blocks_2_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_2_add_1 signals
// --------------------------
logic [stream_blocks_2_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_2_add_1_mdata_in_0        [stream_blocks_2_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_2_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_2_add_1_edata_in_0;
logic                             stream_blocks_2_add_1_data_in_0_valid;
logic                             stream_blocks_2_add_1_data_in_0_ready;
logic [stream_blocks_2_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_2_add_1_mdata_in_1        [stream_blocks_2_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_2_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_2_add_1_edata_in_1;
logic                             stream_blocks_2_add_1_data_in_1_valid;
logic                             stream_blocks_2_add_1_data_in_1_ready;
logic [stream_blocks_2_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_2_add_1_mdata_out_0        [stream_blocks_2_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_2_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_2_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_2_add_1_edata_out_0;
logic                             stream_blocks_2_add_1_data_out_0_valid;
logic                             stream_blocks_2_add_1_data_out_0_ready;
// --------------------------
//   fork2_6 signals
// --------------------------
logic [fork2_6_DATA_IN_0_PRECISION_0-1:0]  fork2_6_mdata_in_0        [fork2_6_DATA_IN_0_PARALLELISM_DIM_0*fork2_6_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_6_DATA_IN_0_PRECISION_1-1:0]  fork2_6_edata_in_0;
logic                             fork2_6_data_in_0_valid;
logic                             fork2_6_data_in_0_ready;
logic [fork2_6_DATA_OUT_0_PRECISION_0-1:0]  fork2_6_mdata_out_0        [fork2_6_DATA_OUT_0_PARALLELISM_DIM_0*fork2_6_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_6_DATA_OUT_0_PRECISION_1-1:0]  fork2_6_edata_out_0;
logic                             fork2_6_data_out_0_valid;
logic                             fork2_6_data_out_0_ready;
logic [fork2_6_DATA_OUT_1_PRECISION_0-1:0]  fork2_6_mdata_out_1        [fork2_6_DATA_OUT_1_PARALLELISM_DIM_0*fork2_6_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_6_DATA_OUT_1_PRECISION_1-1:0]  fork2_6_edata_out_1;
logic                             fork2_6_data_out_1_valid;
logic                             fork2_6_data_out_1_ready;
// --------------------------
//   stream_blocks_3_linear1 signals
// --------------------------
logic [stream_blocks_3_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_3_linear1_mdata_in_0        [stream_blocks_3_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_3_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_3_linear1_edata_in_0;
logic                             stream_blocks_3_linear1_data_in_0_valid;
logic                             stream_blocks_3_linear1_data_in_0_ready;
logic [stream_blocks_3_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_3_linear1_mweight        [stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_3_linear1_eweight;
logic                             stream_blocks_3_linear1_weight_valid;
logic                             stream_blocks_3_linear1_weight_ready;
logic [stream_blocks_3_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_3_linear1_mbias        [stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_3_linear1_ebias;
logic                             stream_blocks_3_linear1_bias_valid;
logic                             stream_blocks_3_linear1_bias_ready;
logic [stream_blocks_3_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_3_linear1_mdata_out_0        [stream_blocks_3_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_3_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_3_linear1_edata_out_0;
logic                             stream_blocks_3_linear1_data_out_0_valid;
logic                             stream_blocks_3_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_3_act signals
// --------------------------
logic [stream_blocks_3_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_3_act_mdata_in_0        [stream_blocks_3_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_3_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_3_act_edata_in_0;
logic                             stream_blocks_3_act_data_in_0_valid;
logic                             stream_blocks_3_act_data_in_0_ready;
logic [stream_blocks_3_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_3_act_mdata_out_0        [stream_blocks_3_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_3_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_3_act_edata_out_0;
logic                             stream_blocks_3_act_data_out_0_valid;
logic                             stream_blocks_3_act_data_out_0_ready;
// --------------------------
//   stream_blocks_3_linear2 signals
// --------------------------
logic [stream_blocks_3_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_3_linear2_mdata_in_0        [stream_blocks_3_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_3_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_3_linear2_edata_in_0;
logic                             stream_blocks_3_linear2_data_in_0_valid;
logic                             stream_blocks_3_linear2_data_in_0_ready;
logic [stream_blocks_3_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_3_linear2_mweight        [stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_3_linear2_eweight;
logic                             stream_blocks_3_linear2_weight_valid;
logic                             stream_blocks_3_linear2_weight_ready;
logic [stream_blocks_3_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_3_linear2_mbias        [stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_3_linear2_ebias;
logic                             stream_blocks_3_linear2_bias_valid;
logic                             stream_blocks_3_linear2_bias_ready;
logic [stream_blocks_3_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_3_linear2_mdata_out_0        [stream_blocks_3_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_3_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_3_linear2_edata_out_0;
logic                             stream_blocks_3_linear2_data_out_0_valid;
logic                             stream_blocks_3_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_3_norm1 signals
// --------------------------
logic [stream_blocks_3_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_3_norm1_mdata_in_0        [stream_blocks_3_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_3_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_3_norm1_edata_in_0;
logic                             stream_blocks_3_norm1_data_in_0_valid;
logic                             stream_blocks_3_norm1_data_in_0_ready;
logic [stream_blocks_3_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_3_norm1_mweight        [stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_3_norm1_eweight;
logic                             stream_blocks_3_norm1_weight_valid;
logic                             stream_blocks_3_norm1_weight_ready;
logic [stream_blocks_3_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_3_norm1_mbias        [stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_3_norm1_ebias;
logic                             stream_blocks_3_norm1_bias_valid;
logic                             stream_blocks_3_norm1_bias_ready;
logic [stream_blocks_3_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_3_norm1_mdata_out_0        [stream_blocks_3_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_3_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_3_norm1_edata_out_0;
logic                             stream_blocks_3_norm1_data_out_0_valid;
logic                             stream_blocks_3_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_3_add signals
// --------------------------
logic [stream_blocks_3_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_3_add_mdata_in_0        [stream_blocks_3_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_3_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_3_add_edata_in_0;
logic                             stream_blocks_3_add_data_in_0_valid;
logic                             stream_blocks_3_add_data_in_0_ready;
logic [stream_blocks_3_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_3_add_mdata_in_1        [stream_blocks_3_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_3_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_3_add_edata_in_1;
logic                             stream_blocks_3_add_data_in_1_valid;
logic                             stream_blocks_3_add_data_in_1_ready;
logic [stream_blocks_3_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_3_add_mdata_out_0        [stream_blocks_3_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_3_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_3_add_edata_out_0;
logic                             stream_blocks_3_add_data_out_0_valid;
logic                             stream_blocks_3_add_data_out_0_ready;
// --------------------------
//   fork2_7 signals
// --------------------------
logic [fork2_7_DATA_IN_0_PRECISION_0-1:0]  fork2_7_mdata_in_0        [fork2_7_DATA_IN_0_PARALLELISM_DIM_0*fork2_7_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_7_DATA_IN_0_PRECISION_1-1:0]  fork2_7_edata_in_0;
logic                             fork2_7_data_in_0_valid;
logic                             fork2_7_data_in_0_ready;
logic [fork2_7_DATA_OUT_0_PRECISION_0-1:0]  fork2_7_mdata_out_0        [fork2_7_DATA_OUT_0_PARALLELISM_DIM_0*fork2_7_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_7_DATA_OUT_0_PRECISION_1-1:0]  fork2_7_edata_out_0;
logic                             fork2_7_data_out_0_valid;
logic                             fork2_7_data_out_0_ready;
logic [fork2_7_DATA_OUT_1_PRECISION_0-1:0]  fork2_7_mdata_out_1        [fork2_7_DATA_OUT_1_PARALLELISM_DIM_0*fork2_7_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_7_DATA_OUT_1_PRECISION_1-1:0]  fork2_7_edata_out_1;
logic                             fork2_7_data_out_1_valid;
logic                             fork2_7_data_out_1_ready;
// --------------------------
//   stream_blocks_3_attention signals
// --------------------------
logic [stream_blocks_3_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_3_attention_mdata_in_0        [stream_blocks_3_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_3_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_3_attention_edata_in_0;
logic                             stream_blocks_3_attention_data_in_0_valid;
logic                             stream_blocks_3_attention_data_in_0_ready;
logic [stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_3_attention_mquery_weight        [stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_3_attention_equery_weight;
logic                             stream_blocks_3_attention_query_weight_valid;
logic                             stream_blocks_3_attention_query_weight_ready;
logic [stream_blocks_3_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_3_attention_mquery_bias        [stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_3_attention_equery_bias;
logic                             stream_blocks_3_attention_query_bias_valid;
logic                             stream_blocks_3_attention_query_bias_ready;
logic [stream_blocks_3_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_3_attention_mkey_weight        [stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_3_attention_ekey_weight;
logic                             stream_blocks_3_attention_key_weight_valid;
logic                             stream_blocks_3_attention_key_weight_ready;
logic [stream_blocks_3_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_3_attention_mkey_bias        [stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_3_attention_ekey_bias;
logic                             stream_blocks_3_attention_key_bias_valid;
logic                             stream_blocks_3_attention_key_bias_ready;
logic [stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_3_attention_mvalue_weight        [stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_3_attention_evalue_weight;
logic                             stream_blocks_3_attention_value_weight_valid;
logic                             stream_blocks_3_attention_value_weight_ready;
logic [stream_blocks_3_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_3_attention_mvalue_bias        [stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_3_attention_evalue_bias;
logic                             stream_blocks_3_attention_value_bias_valid;
logic                             stream_blocks_3_attention_value_bias_ready;
logic [stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_3_attention_mproj_weight        [stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_3_attention_eproj_weight;
logic                             stream_blocks_3_attention_proj_weight_valid;
logic                             stream_blocks_3_attention_proj_weight_ready;
logic [stream_blocks_3_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_3_attention_mproj_bias        [stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_3_attention_eproj_bias;
logic                             stream_blocks_3_attention_proj_bias_valid;
logic                             stream_blocks_3_attention_proj_bias_ready;
logic [stream_blocks_3_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_3_attention_mdata_out_0        [stream_blocks_3_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_3_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_3_attention_edata_out_0;
logic                             stream_blocks_3_attention_data_out_0_valid;
logic                             stream_blocks_3_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_3_norm2 signals
// --------------------------
logic [stream_blocks_3_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_3_norm2_mdata_in_0        [stream_blocks_3_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_3_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_3_norm2_edata_in_0;
logic                             stream_blocks_3_norm2_data_in_0_valid;
logic                             stream_blocks_3_norm2_data_in_0_ready;
logic [stream_blocks_3_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_3_norm2_mweight        [stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_3_norm2_eweight;
logic                             stream_blocks_3_norm2_weight_valid;
logic                             stream_blocks_3_norm2_weight_ready;
logic [stream_blocks_3_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_3_norm2_mbias        [stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_3_norm2_ebias;
logic                             stream_blocks_3_norm2_bias_valid;
logic                             stream_blocks_3_norm2_bias_ready;
logic [stream_blocks_3_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_3_norm2_mdata_out_0        [stream_blocks_3_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_3_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_3_norm2_edata_out_0;
logic                             stream_blocks_3_norm2_data_out_0_valid;
logic                             stream_blocks_3_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_3_add_1 signals
// --------------------------
logic [stream_blocks_3_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_3_add_1_mdata_in_0        [stream_blocks_3_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_3_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_3_add_1_edata_in_0;
logic                             stream_blocks_3_add_1_data_in_0_valid;
logic                             stream_blocks_3_add_1_data_in_0_ready;
logic [stream_blocks_3_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_3_add_1_mdata_in_1        [stream_blocks_3_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_3_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_3_add_1_edata_in_1;
logic                             stream_blocks_3_add_1_data_in_1_valid;
logic                             stream_blocks_3_add_1_data_in_1_ready;
logic [stream_blocks_3_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_3_add_1_mdata_out_0        [stream_blocks_3_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_3_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_3_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_3_add_1_edata_out_0;
logic                             stream_blocks_3_add_1_data_out_0_valid;
logic                             stream_blocks_3_add_1_data_out_0_ready;
// --------------------------
//   fork2_8 signals
// --------------------------
logic [fork2_8_DATA_IN_0_PRECISION_0-1:0]  fork2_8_mdata_in_0        [fork2_8_DATA_IN_0_PARALLELISM_DIM_0*fork2_8_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_8_DATA_IN_0_PRECISION_1-1:0]  fork2_8_edata_in_0;
logic                             fork2_8_data_in_0_valid;
logic                             fork2_8_data_in_0_ready;
logic [fork2_8_DATA_OUT_0_PRECISION_0-1:0]  fork2_8_mdata_out_0        [fork2_8_DATA_OUT_0_PARALLELISM_DIM_0*fork2_8_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_8_DATA_OUT_0_PRECISION_1-1:0]  fork2_8_edata_out_0;
logic                             fork2_8_data_out_0_valid;
logic                             fork2_8_data_out_0_ready;
logic [fork2_8_DATA_OUT_1_PRECISION_0-1:0]  fork2_8_mdata_out_1        [fork2_8_DATA_OUT_1_PARALLELISM_DIM_0*fork2_8_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_8_DATA_OUT_1_PRECISION_1-1:0]  fork2_8_edata_out_1;
logic                             fork2_8_data_out_1_valid;
logic                             fork2_8_data_out_1_ready;
// --------------------------
//   stream_blocks_4_linear1 signals
// --------------------------
logic [stream_blocks_4_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_4_linear1_mdata_in_0        [stream_blocks_4_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_4_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_4_linear1_edata_in_0;
logic                             stream_blocks_4_linear1_data_in_0_valid;
logic                             stream_blocks_4_linear1_data_in_0_ready;
logic [stream_blocks_4_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_4_linear1_mweight        [stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_4_linear1_eweight;
logic                             stream_blocks_4_linear1_weight_valid;
logic                             stream_blocks_4_linear1_weight_ready;
logic [stream_blocks_4_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_4_linear1_mbias        [stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_4_linear1_ebias;
logic                             stream_blocks_4_linear1_bias_valid;
logic                             stream_blocks_4_linear1_bias_ready;
logic [stream_blocks_4_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_4_linear1_mdata_out_0        [stream_blocks_4_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_4_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_4_linear1_edata_out_0;
logic                             stream_blocks_4_linear1_data_out_0_valid;
logic                             stream_blocks_4_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_4_act signals
// --------------------------
logic [stream_blocks_4_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_4_act_mdata_in_0        [stream_blocks_4_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_4_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_4_act_edata_in_0;
logic                             stream_blocks_4_act_data_in_0_valid;
logic                             stream_blocks_4_act_data_in_0_ready;
logic [stream_blocks_4_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_4_act_mdata_out_0        [stream_blocks_4_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_4_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_4_act_edata_out_0;
logic                             stream_blocks_4_act_data_out_0_valid;
logic                             stream_blocks_4_act_data_out_0_ready;
// --------------------------
//   stream_blocks_4_linear2 signals
// --------------------------
logic [stream_blocks_4_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_4_linear2_mdata_in_0        [stream_blocks_4_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_4_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_4_linear2_edata_in_0;
logic                             stream_blocks_4_linear2_data_in_0_valid;
logic                             stream_blocks_4_linear2_data_in_0_ready;
logic [stream_blocks_4_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_4_linear2_mweight        [stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_4_linear2_eweight;
logic                             stream_blocks_4_linear2_weight_valid;
logic                             stream_blocks_4_linear2_weight_ready;
logic [stream_blocks_4_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_4_linear2_mbias        [stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_4_linear2_ebias;
logic                             stream_blocks_4_linear2_bias_valid;
logic                             stream_blocks_4_linear2_bias_ready;
logic [stream_blocks_4_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_4_linear2_mdata_out_0        [stream_blocks_4_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_4_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_4_linear2_edata_out_0;
logic                             stream_blocks_4_linear2_data_out_0_valid;
logic                             stream_blocks_4_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_4_norm1 signals
// --------------------------
logic [stream_blocks_4_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_4_norm1_mdata_in_0        [stream_blocks_4_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_4_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_4_norm1_edata_in_0;
logic                             stream_blocks_4_norm1_data_in_0_valid;
logic                             stream_blocks_4_norm1_data_in_0_ready;
logic [stream_blocks_4_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_4_norm1_mweight        [stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_4_norm1_eweight;
logic                             stream_blocks_4_norm1_weight_valid;
logic                             stream_blocks_4_norm1_weight_ready;
logic [stream_blocks_4_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_4_norm1_mbias        [stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_4_norm1_ebias;
logic                             stream_blocks_4_norm1_bias_valid;
logic                             stream_blocks_4_norm1_bias_ready;
logic [stream_blocks_4_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_4_norm1_mdata_out_0        [stream_blocks_4_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_4_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_4_norm1_edata_out_0;
logic                             stream_blocks_4_norm1_data_out_0_valid;
logic                             stream_blocks_4_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_4_add signals
// --------------------------
logic [stream_blocks_4_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_4_add_mdata_in_0        [stream_blocks_4_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_4_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_4_add_edata_in_0;
logic                             stream_blocks_4_add_data_in_0_valid;
logic                             stream_blocks_4_add_data_in_0_ready;
logic [stream_blocks_4_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_4_add_mdata_in_1        [stream_blocks_4_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_4_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_4_add_edata_in_1;
logic                             stream_blocks_4_add_data_in_1_valid;
logic                             stream_blocks_4_add_data_in_1_ready;
logic [stream_blocks_4_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_4_add_mdata_out_0        [stream_blocks_4_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_4_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_4_add_edata_out_0;
logic                             stream_blocks_4_add_data_out_0_valid;
logic                             stream_blocks_4_add_data_out_0_ready;
// --------------------------
//   fork2_9 signals
// --------------------------
logic [fork2_9_DATA_IN_0_PRECISION_0-1:0]  fork2_9_mdata_in_0        [fork2_9_DATA_IN_0_PARALLELISM_DIM_0*fork2_9_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_9_DATA_IN_0_PRECISION_1-1:0]  fork2_9_edata_in_0;
logic                             fork2_9_data_in_0_valid;
logic                             fork2_9_data_in_0_ready;
logic [fork2_9_DATA_OUT_0_PRECISION_0-1:0]  fork2_9_mdata_out_0        [fork2_9_DATA_OUT_0_PARALLELISM_DIM_0*fork2_9_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_9_DATA_OUT_0_PRECISION_1-1:0]  fork2_9_edata_out_0;
logic                             fork2_9_data_out_0_valid;
logic                             fork2_9_data_out_0_ready;
logic [fork2_9_DATA_OUT_1_PRECISION_0-1:0]  fork2_9_mdata_out_1        [fork2_9_DATA_OUT_1_PARALLELISM_DIM_0*fork2_9_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_9_DATA_OUT_1_PRECISION_1-1:0]  fork2_9_edata_out_1;
logic                             fork2_9_data_out_1_valid;
logic                             fork2_9_data_out_1_ready;
// --------------------------
//   stream_blocks_4_attention signals
// --------------------------
logic [stream_blocks_4_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_4_attention_mdata_in_0        [stream_blocks_4_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_4_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_4_attention_edata_in_0;
logic                             stream_blocks_4_attention_data_in_0_valid;
logic                             stream_blocks_4_attention_data_in_0_ready;
logic [stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_4_attention_mquery_weight        [stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_4_attention_equery_weight;
logic                             stream_blocks_4_attention_query_weight_valid;
logic                             stream_blocks_4_attention_query_weight_ready;
logic [stream_blocks_4_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_4_attention_mquery_bias        [stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_4_attention_equery_bias;
logic                             stream_blocks_4_attention_query_bias_valid;
logic                             stream_blocks_4_attention_query_bias_ready;
logic [stream_blocks_4_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_4_attention_mkey_weight        [stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_4_attention_ekey_weight;
logic                             stream_blocks_4_attention_key_weight_valid;
logic                             stream_blocks_4_attention_key_weight_ready;
logic [stream_blocks_4_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_4_attention_mkey_bias        [stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_4_attention_ekey_bias;
logic                             stream_blocks_4_attention_key_bias_valid;
logic                             stream_blocks_4_attention_key_bias_ready;
logic [stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_4_attention_mvalue_weight        [stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_4_attention_evalue_weight;
logic                             stream_blocks_4_attention_value_weight_valid;
logic                             stream_blocks_4_attention_value_weight_ready;
logic [stream_blocks_4_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_4_attention_mvalue_bias        [stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_4_attention_evalue_bias;
logic                             stream_blocks_4_attention_value_bias_valid;
logic                             stream_blocks_4_attention_value_bias_ready;
logic [stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_4_attention_mproj_weight        [stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_4_attention_eproj_weight;
logic                             stream_blocks_4_attention_proj_weight_valid;
logic                             stream_blocks_4_attention_proj_weight_ready;
logic [stream_blocks_4_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_4_attention_mproj_bias        [stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_4_attention_eproj_bias;
logic                             stream_blocks_4_attention_proj_bias_valid;
logic                             stream_blocks_4_attention_proj_bias_ready;
logic [stream_blocks_4_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_4_attention_mdata_out_0        [stream_blocks_4_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_4_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_4_attention_edata_out_0;
logic                             stream_blocks_4_attention_data_out_0_valid;
logic                             stream_blocks_4_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_4_norm2 signals
// --------------------------
logic [stream_blocks_4_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_4_norm2_mdata_in_0        [stream_blocks_4_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_4_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_4_norm2_edata_in_0;
logic                             stream_blocks_4_norm2_data_in_0_valid;
logic                             stream_blocks_4_norm2_data_in_0_ready;
logic [stream_blocks_4_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_4_norm2_mweight        [stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_4_norm2_eweight;
logic                             stream_blocks_4_norm2_weight_valid;
logic                             stream_blocks_4_norm2_weight_ready;
logic [stream_blocks_4_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_4_norm2_mbias        [stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_4_norm2_ebias;
logic                             stream_blocks_4_norm2_bias_valid;
logic                             stream_blocks_4_norm2_bias_ready;
logic [stream_blocks_4_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_4_norm2_mdata_out_0        [stream_blocks_4_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_4_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_4_norm2_edata_out_0;
logic                             stream_blocks_4_norm2_data_out_0_valid;
logic                             stream_blocks_4_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_4_add_1 signals
// --------------------------
logic [stream_blocks_4_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_4_add_1_mdata_in_0        [stream_blocks_4_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_4_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_4_add_1_edata_in_0;
logic                             stream_blocks_4_add_1_data_in_0_valid;
logic                             stream_blocks_4_add_1_data_in_0_ready;
logic [stream_blocks_4_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_4_add_1_mdata_in_1        [stream_blocks_4_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_4_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_4_add_1_edata_in_1;
logic                             stream_blocks_4_add_1_data_in_1_valid;
logic                             stream_blocks_4_add_1_data_in_1_ready;
logic [stream_blocks_4_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_4_add_1_mdata_out_0        [stream_blocks_4_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_4_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_4_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_4_add_1_edata_out_0;
logic                             stream_blocks_4_add_1_data_out_0_valid;
logic                             stream_blocks_4_add_1_data_out_0_ready;
// --------------------------
//   fork2_10 signals
// --------------------------
logic [fork2_10_DATA_IN_0_PRECISION_0-1:0]  fork2_10_mdata_in_0        [fork2_10_DATA_IN_0_PARALLELISM_DIM_0*fork2_10_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_10_DATA_IN_0_PRECISION_1-1:0]  fork2_10_edata_in_0;
logic                             fork2_10_data_in_0_valid;
logic                             fork2_10_data_in_0_ready;
logic [fork2_10_DATA_OUT_0_PRECISION_0-1:0]  fork2_10_mdata_out_0        [fork2_10_DATA_OUT_0_PARALLELISM_DIM_0*fork2_10_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_10_DATA_OUT_0_PRECISION_1-1:0]  fork2_10_edata_out_0;
logic                             fork2_10_data_out_0_valid;
logic                             fork2_10_data_out_0_ready;
logic [fork2_10_DATA_OUT_1_PRECISION_0-1:0]  fork2_10_mdata_out_1        [fork2_10_DATA_OUT_1_PARALLELISM_DIM_0*fork2_10_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_10_DATA_OUT_1_PRECISION_1-1:0]  fork2_10_edata_out_1;
logic                             fork2_10_data_out_1_valid;
logic                             fork2_10_data_out_1_ready;
// --------------------------
//   stream_blocks_5_linear1 signals
// --------------------------
logic [stream_blocks_5_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_5_linear1_mdata_in_0        [stream_blocks_5_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_5_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_5_linear1_edata_in_0;
logic                             stream_blocks_5_linear1_data_in_0_valid;
logic                             stream_blocks_5_linear1_data_in_0_ready;
logic [stream_blocks_5_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_5_linear1_mweight        [stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_5_linear1_eweight;
logic                             stream_blocks_5_linear1_weight_valid;
logic                             stream_blocks_5_linear1_weight_ready;
logic [stream_blocks_5_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_5_linear1_mbias        [stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_5_linear1_ebias;
logic                             stream_blocks_5_linear1_bias_valid;
logic                             stream_blocks_5_linear1_bias_ready;
logic [stream_blocks_5_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_5_linear1_mdata_out_0        [stream_blocks_5_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_5_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_5_linear1_edata_out_0;
logic                             stream_blocks_5_linear1_data_out_0_valid;
logic                             stream_blocks_5_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_5_act signals
// --------------------------
logic [stream_blocks_5_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_5_act_mdata_in_0        [stream_blocks_5_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_5_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_5_act_edata_in_0;
logic                             stream_blocks_5_act_data_in_0_valid;
logic                             stream_blocks_5_act_data_in_0_ready;
logic [stream_blocks_5_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_5_act_mdata_out_0        [stream_blocks_5_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_5_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_5_act_edata_out_0;
logic                             stream_blocks_5_act_data_out_0_valid;
logic                             stream_blocks_5_act_data_out_0_ready;
// --------------------------
//   stream_blocks_5_linear2 signals
// --------------------------
logic [stream_blocks_5_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_5_linear2_mdata_in_0        [stream_blocks_5_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_5_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_5_linear2_edata_in_0;
logic                             stream_blocks_5_linear2_data_in_0_valid;
logic                             stream_blocks_5_linear2_data_in_0_ready;
logic [stream_blocks_5_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_5_linear2_mweight        [stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_5_linear2_eweight;
logic                             stream_blocks_5_linear2_weight_valid;
logic                             stream_blocks_5_linear2_weight_ready;
logic [stream_blocks_5_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_5_linear2_mbias        [stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_5_linear2_ebias;
logic                             stream_blocks_5_linear2_bias_valid;
logic                             stream_blocks_5_linear2_bias_ready;
logic [stream_blocks_5_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_5_linear2_mdata_out_0        [stream_blocks_5_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_5_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_5_linear2_edata_out_0;
logic                             stream_blocks_5_linear2_data_out_0_valid;
logic                             stream_blocks_5_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_5_norm1 signals
// --------------------------
logic [stream_blocks_5_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_5_norm1_mdata_in_0        [stream_blocks_5_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_5_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_5_norm1_edata_in_0;
logic                             stream_blocks_5_norm1_data_in_0_valid;
logic                             stream_blocks_5_norm1_data_in_0_ready;
logic [stream_blocks_5_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_5_norm1_mweight        [stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_5_norm1_eweight;
logic                             stream_blocks_5_norm1_weight_valid;
logic                             stream_blocks_5_norm1_weight_ready;
logic [stream_blocks_5_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_5_norm1_mbias        [stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_5_norm1_ebias;
logic                             stream_blocks_5_norm1_bias_valid;
logic                             stream_blocks_5_norm1_bias_ready;
logic [stream_blocks_5_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_5_norm1_mdata_out_0        [stream_blocks_5_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_5_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_5_norm1_edata_out_0;
logic                             stream_blocks_5_norm1_data_out_0_valid;
logic                             stream_blocks_5_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_5_add signals
// --------------------------
logic [stream_blocks_5_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_5_add_mdata_in_0        [stream_blocks_5_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_5_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_5_add_edata_in_0;
logic                             stream_blocks_5_add_data_in_0_valid;
logic                             stream_blocks_5_add_data_in_0_ready;
logic [stream_blocks_5_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_5_add_mdata_in_1        [stream_blocks_5_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_5_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_5_add_edata_in_1;
logic                             stream_blocks_5_add_data_in_1_valid;
logic                             stream_blocks_5_add_data_in_1_ready;
logic [stream_blocks_5_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_5_add_mdata_out_0        [stream_blocks_5_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_5_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_5_add_edata_out_0;
logic                             stream_blocks_5_add_data_out_0_valid;
logic                             stream_blocks_5_add_data_out_0_ready;
// --------------------------
//   fork2_11 signals
// --------------------------
logic [fork2_11_DATA_IN_0_PRECISION_0-1:0]  fork2_11_mdata_in_0        [fork2_11_DATA_IN_0_PARALLELISM_DIM_0*fork2_11_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_11_DATA_IN_0_PRECISION_1-1:0]  fork2_11_edata_in_0;
logic                             fork2_11_data_in_0_valid;
logic                             fork2_11_data_in_0_ready;
logic [fork2_11_DATA_OUT_0_PRECISION_0-1:0]  fork2_11_mdata_out_0        [fork2_11_DATA_OUT_0_PARALLELISM_DIM_0*fork2_11_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_11_DATA_OUT_0_PRECISION_1-1:0]  fork2_11_edata_out_0;
logic                             fork2_11_data_out_0_valid;
logic                             fork2_11_data_out_0_ready;
logic [fork2_11_DATA_OUT_1_PRECISION_0-1:0]  fork2_11_mdata_out_1        [fork2_11_DATA_OUT_1_PARALLELISM_DIM_0*fork2_11_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_11_DATA_OUT_1_PRECISION_1-1:0]  fork2_11_edata_out_1;
logic                             fork2_11_data_out_1_valid;
logic                             fork2_11_data_out_1_ready;
// --------------------------
//   stream_blocks_5_attention signals
// --------------------------
logic [stream_blocks_5_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_5_attention_mdata_in_0        [stream_blocks_5_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_5_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_5_attention_edata_in_0;
logic                             stream_blocks_5_attention_data_in_0_valid;
logic                             stream_blocks_5_attention_data_in_0_ready;
logic [stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_5_attention_mquery_weight        [stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_5_attention_equery_weight;
logic                             stream_blocks_5_attention_query_weight_valid;
logic                             stream_blocks_5_attention_query_weight_ready;
logic [stream_blocks_5_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_5_attention_mquery_bias        [stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_5_attention_equery_bias;
logic                             stream_blocks_5_attention_query_bias_valid;
logic                             stream_blocks_5_attention_query_bias_ready;
logic [stream_blocks_5_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_5_attention_mkey_weight        [stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_5_attention_ekey_weight;
logic                             stream_blocks_5_attention_key_weight_valid;
logic                             stream_blocks_5_attention_key_weight_ready;
logic [stream_blocks_5_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_5_attention_mkey_bias        [stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_5_attention_ekey_bias;
logic                             stream_blocks_5_attention_key_bias_valid;
logic                             stream_blocks_5_attention_key_bias_ready;
logic [stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_5_attention_mvalue_weight        [stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_5_attention_evalue_weight;
logic                             stream_blocks_5_attention_value_weight_valid;
logic                             stream_blocks_5_attention_value_weight_ready;
logic [stream_blocks_5_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_5_attention_mvalue_bias        [stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_5_attention_evalue_bias;
logic                             stream_blocks_5_attention_value_bias_valid;
logic                             stream_blocks_5_attention_value_bias_ready;
logic [stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_5_attention_mproj_weight        [stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_5_attention_eproj_weight;
logic                             stream_blocks_5_attention_proj_weight_valid;
logic                             stream_blocks_5_attention_proj_weight_ready;
logic [stream_blocks_5_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_5_attention_mproj_bias        [stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_5_attention_eproj_bias;
logic                             stream_blocks_5_attention_proj_bias_valid;
logic                             stream_blocks_5_attention_proj_bias_ready;
logic [stream_blocks_5_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_5_attention_mdata_out_0        [stream_blocks_5_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_5_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_5_attention_edata_out_0;
logic                             stream_blocks_5_attention_data_out_0_valid;
logic                             stream_blocks_5_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_5_norm2 signals
// --------------------------
logic [stream_blocks_5_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_5_norm2_mdata_in_0        [stream_blocks_5_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_5_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_5_norm2_edata_in_0;
logic                             stream_blocks_5_norm2_data_in_0_valid;
logic                             stream_blocks_5_norm2_data_in_0_ready;
logic [stream_blocks_5_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_5_norm2_mweight        [stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_5_norm2_eweight;
logic                             stream_blocks_5_norm2_weight_valid;
logic                             stream_blocks_5_norm2_weight_ready;
logic [stream_blocks_5_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_5_norm2_mbias        [stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_5_norm2_ebias;
logic                             stream_blocks_5_norm2_bias_valid;
logic                             stream_blocks_5_norm2_bias_ready;
logic [stream_blocks_5_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_5_norm2_mdata_out_0        [stream_blocks_5_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_5_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_5_norm2_edata_out_0;
logic                             stream_blocks_5_norm2_data_out_0_valid;
logic                             stream_blocks_5_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_5_add_1 signals
// --------------------------
logic [stream_blocks_5_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_5_add_1_mdata_in_0        [stream_blocks_5_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_5_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_5_add_1_edata_in_0;
logic                             stream_blocks_5_add_1_data_in_0_valid;
logic                             stream_blocks_5_add_1_data_in_0_ready;
logic [stream_blocks_5_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_5_add_1_mdata_in_1        [stream_blocks_5_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_5_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_5_add_1_edata_in_1;
logic                             stream_blocks_5_add_1_data_in_1_valid;
logic                             stream_blocks_5_add_1_data_in_1_ready;
logic [stream_blocks_5_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_5_add_1_mdata_out_0        [stream_blocks_5_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_5_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_5_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_5_add_1_edata_out_0;
logic                             stream_blocks_5_add_1_data_out_0_valid;
logic                             stream_blocks_5_add_1_data_out_0_ready;
// --------------------------
//   fork2_12 signals
// --------------------------
logic [fork2_12_DATA_IN_0_PRECISION_0-1:0]  fork2_12_mdata_in_0        [fork2_12_DATA_IN_0_PARALLELISM_DIM_0*fork2_12_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_12_DATA_IN_0_PRECISION_1-1:0]  fork2_12_edata_in_0;
logic                             fork2_12_data_in_0_valid;
logic                             fork2_12_data_in_0_ready;
logic [fork2_12_DATA_OUT_0_PRECISION_0-1:0]  fork2_12_mdata_out_0        [fork2_12_DATA_OUT_0_PARALLELISM_DIM_0*fork2_12_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_12_DATA_OUT_0_PRECISION_1-1:0]  fork2_12_edata_out_0;
logic                             fork2_12_data_out_0_valid;
logic                             fork2_12_data_out_0_ready;
logic [fork2_12_DATA_OUT_1_PRECISION_0-1:0]  fork2_12_mdata_out_1        [fork2_12_DATA_OUT_1_PARALLELISM_DIM_0*fork2_12_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_12_DATA_OUT_1_PRECISION_1-1:0]  fork2_12_edata_out_1;
logic                             fork2_12_data_out_1_valid;
logic                             fork2_12_data_out_1_ready;
// --------------------------
//   stream_blocks_6_linear1 signals
// --------------------------
logic [stream_blocks_6_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_6_linear1_mdata_in_0        [stream_blocks_6_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_6_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_6_linear1_edata_in_0;
logic                             stream_blocks_6_linear1_data_in_0_valid;
logic                             stream_blocks_6_linear1_data_in_0_ready;
logic [stream_blocks_6_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_6_linear1_mweight        [stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_6_linear1_eweight;
logic                             stream_blocks_6_linear1_weight_valid;
logic                             stream_blocks_6_linear1_weight_ready;
logic [stream_blocks_6_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_6_linear1_mbias        [stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_6_linear1_ebias;
logic                             stream_blocks_6_linear1_bias_valid;
logic                             stream_blocks_6_linear1_bias_ready;
logic [stream_blocks_6_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_6_linear1_mdata_out_0        [stream_blocks_6_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_6_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_6_linear1_edata_out_0;
logic                             stream_blocks_6_linear1_data_out_0_valid;
logic                             stream_blocks_6_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_6_act signals
// --------------------------
logic [stream_blocks_6_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_6_act_mdata_in_0        [stream_blocks_6_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_6_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_6_act_edata_in_0;
logic                             stream_blocks_6_act_data_in_0_valid;
logic                             stream_blocks_6_act_data_in_0_ready;
logic [stream_blocks_6_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_6_act_mdata_out_0        [stream_blocks_6_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_6_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_6_act_edata_out_0;
logic                             stream_blocks_6_act_data_out_0_valid;
logic                             stream_blocks_6_act_data_out_0_ready;
// --------------------------
//   stream_blocks_6_linear2 signals
// --------------------------
logic [stream_blocks_6_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_6_linear2_mdata_in_0        [stream_blocks_6_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_6_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_6_linear2_edata_in_0;
logic                             stream_blocks_6_linear2_data_in_0_valid;
logic                             stream_blocks_6_linear2_data_in_0_ready;
logic [stream_blocks_6_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_6_linear2_mweight        [stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_6_linear2_eweight;
logic                             stream_blocks_6_linear2_weight_valid;
logic                             stream_blocks_6_linear2_weight_ready;
logic [stream_blocks_6_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_6_linear2_mbias        [stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_6_linear2_ebias;
logic                             stream_blocks_6_linear2_bias_valid;
logic                             stream_blocks_6_linear2_bias_ready;
logic [stream_blocks_6_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_6_linear2_mdata_out_0        [stream_blocks_6_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_6_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_6_linear2_edata_out_0;
logic                             stream_blocks_6_linear2_data_out_0_valid;
logic                             stream_blocks_6_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_6_norm1 signals
// --------------------------
logic [stream_blocks_6_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_6_norm1_mdata_in_0        [stream_blocks_6_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_6_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_6_norm1_edata_in_0;
logic                             stream_blocks_6_norm1_data_in_0_valid;
logic                             stream_blocks_6_norm1_data_in_0_ready;
logic [stream_blocks_6_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_6_norm1_mweight        [stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_6_norm1_eweight;
logic                             stream_blocks_6_norm1_weight_valid;
logic                             stream_blocks_6_norm1_weight_ready;
logic [stream_blocks_6_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_6_norm1_mbias        [stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_6_norm1_ebias;
logic                             stream_blocks_6_norm1_bias_valid;
logic                             stream_blocks_6_norm1_bias_ready;
logic [stream_blocks_6_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_6_norm1_mdata_out_0        [stream_blocks_6_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_6_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_6_norm1_edata_out_0;
logic                             stream_blocks_6_norm1_data_out_0_valid;
logic                             stream_blocks_6_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_6_add signals
// --------------------------
logic [stream_blocks_6_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_6_add_mdata_in_0        [stream_blocks_6_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_6_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_6_add_edata_in_0;
logic                             stream_blocks_6_add_data_in_0_valid;
logic                             stream_blocks_6_add_data_in_0_ready;
logic [stream_blocks_6_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_6_add_mdata_in_1        [stream_blocks_6_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_6_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_6_add_edata_in_1;
logic                             stream_blocks_6_add_data_in_1_valid;
logic                             stream_blocks_6_add_data_in_1_ready;
logic [stream_blocks_6_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_6_add_mdata_out_0        [stream_blocks_6_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_6_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_6_add_edata_out_0;
logic                             stream_blocks_6_add_data_out_0_valid;
logic                             stream_blocks_6_add_data_out_0_ready;
// --------------------------
//   fork2_13 signals
// --------------------------
logic [fork2_13_DATA_IN_0_PRECISION_0-1:0]  fork2_13_mdata_in_0        [fork2_13_DATA_IN_0_PARALLELISM_DIM_0*fork2_13_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_13_DATA_IN_0_PRECISION_1-1:0]  fork2_13_edata_in_0;
logic                             fork2_13_data_in_0_valid;
logic                             fork2_13_data_in_0_ready;
logic [fork2_13_DATA_OUT_0_PRECISION_0-1:0]  fork2_13_mdata_out_0        [fork2_13_DATA_OUT_0_PARALLELISM_DIM_0*fork2_13_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_13_DATA_OUT_0_PRECISION_1-1:0]  fork2_13_edata_out_0;
logic                             fork2_13_data_out_0_valid;
logic                             fork2_13_data_out_0_ready;
logic [fork2_13_DATA_OUT_1_PRECISION_0-1:0]  fork2_13_mdata_out_1        [fork2_13_DATA_OUT_1_PARALLELISM_DIM_0*fork2_13_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_13_DATA_OUT_1_PRECISION_1-1:0]  fork2_13_edata_out_1;
logic                             fork2_13_data_out_1_valid;
logic                             fork2_13_data_out_1_ready;
// --------------------------
//   stream_blocks_6_attention signals
// --------------------------
logic [stream_blocks_6_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_6_attention_mdata_in_0        [stream_blocks_6_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_6_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_6_attention_edata_in_0;
logic                             stream_blocks_6_attention_data_in_0_valid;
logic                             stream_blocks_6_attention_data_in_0_ready;
logic [stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_6_attention_mquery_weight        [stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_6_attention_equery_weight;
logic                             stream_blocks_6_attention_query_weight_valid;
logic                             stream_blocks_6_attention_query_weight_ready;
logic [stream_blocks_6_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_6_attention_mquery_bias        [stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_6_attention_equery_bias;
logic                             stream_blocks_6_attention_query_bias_valid;
logic                             stream_blocks_6_attention_query_bias_ready;
logic [stream_blocks_6_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_6_attention_mkey_weight        [stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_6_attention_ekey_weight;
logic                             stream_blocks_6_attention_key_weight_valid;
logic                             stream_blocks_6_attention_key_weight_ready;
logic [stream_blocks_6_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_6_attention_mkey_bias        [stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_6_attention_ekey_bias;
logic                             stream_blocks_6_attention_key_bias_valid;
logic                             stream_blocks_6_attention_key_bias_ready;
logic [stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_6_attention_mvalue_weight        [stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_6_attention_evalue_weight;
logic                             stream_blocks_6_attention_value_weight_valid;
logic                             stream_blocks_6_attention_value_weight_ready;
logic [stream_blocks_6_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_6_attention_mvalue_bias        [stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_6_attention_evalue_bias;
logic                             stream_blocks_6_attention_value_bias_valid;
logic                             stream_blocks_6_attention_value_bias_ready;
logic [stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_6_attention_mproj_weight        [stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_6_attention_eproj_weight;
logic                             stream_blocks_6_attention_proj_weight_valid;
logic                             stream_blocks_6_attention_proj_weight_ready;
logic [stream_blocks_6_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_6_attention_mproj_bias        [stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_6_attention_eproj_bias;
logic                             stream_blocks_6_attention_proj_bias_valid;
logic                             stream_blocks_6_attention_proj_bias_ready;
logic [stream_blocks_6_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_6_attention_mdata_out_0        [stream_blocks_6_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_6_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_6_attention_edata_out_0;
logic                             stream_blocks_6_attention_data_out_0_valid;
logic                             stream_blocks_6_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_6_norm2 signals
// --------------------------
logic [stream_blocks_6_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_6_norm2_mdata_in_0        [stream_blocks_6_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_6_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_6_norm2_edata_in_0;
logic                             stream_blocks_6_norm2_data_in_0_valid;
logic                             stream_blocks_6_norm2_data_in_0_ready;
logic [stream_blocks_6_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_6_norm2_mweight        [stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_6_norm2_eweight;
logic                             stream_blocks_6_norm2_weight_valid;
logic                             stream_blocks_6_norm2_weight_ready;
logic [stream_blocks_6_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_6_norm2_mbias        [stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_6_norm2_ebias;
logic                             stream_blocks_6_norm2_bias_valid;
logic                             stream_blocks_6_norm2_bias_ready;
logic [stream_blocks_6_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_6_norm2_mdata_out_0        [stream_blocks_6_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_6_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_6_norm2_edata_out_0;
logic                             stream_blocks_6_norm2_data_out_0_valid;
logic                             stream_blocks_6_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_6_add_1 signals
// --------------------------
logic [stream_blocks_6_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_6_add_1_mdata_in_0        [stream_blocks_6_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_6_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_6_add_1_edata_in_0;
logic                             stream_blocks_6_add_1_data_in_0_valid;
logic                             stream_blocks_6_add_1_data_in_0_ready;
logic [stream_blocks_6_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_6_add_1_mdata_in_1        [stream_blocks_6_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_6_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_6_add_1_edata_in_1;
logic                             stream_blocks_6_add_1_data_in_1_valid;
logic                             stream_blocks_6_add_1_data_in_1_ready;
logic [stream_blocks_6_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_6_add_1_mdata_out_0        [stream_blocks_6_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_6_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_6_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_6_add_1_edata_out_0;
logic                             stream_blocks_6_add_1_data_out_0_valid;
logic                             stream_blocks_6_add_1_data_out_0_ready;
// --------------------------
//   fork2_14 signals
// --------------------------
logic [fork2_14_DATA_IN_0_PRECISION_0-1:0]  fork2_14_mdata_in_0        [fork2_14_DATA_IN_0_PARALLELISM_DIM_0*fork2_14_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_14_DATA_IN_0_PRECISION_1-1:0]  fork2_14_edata_in_0;
logic                             fork2_14_data_in_0_valid;
logic                             fork2_14_data_in_0_ready;
logic [fork2_14_DATA_OUT_0_PRECISION_0-1:0]  fork2_14_mdata_out_0        [fork2_14_DATA_OUT_0_PARALLELISM_DIM_0*fork2_14_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_14_DATA_OUT_0_PRECISION_1-1:0]  fork2_14_edata_out_0;
logic                             fork2_14_data_out_0_valid;
logic                             fork2_14_data_out_0_ready;
logic [fork2_14_DATA_OUT_1_PRECISION_0-1:0]  fork2_14_mdata_out_1        [fork2_14_DATA_OUT_1_PARALLELISM_DIM_0*fork2_14_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_14_DATA_OUT_1_PRECISION_1-1:0]  fork2_14_edata_out_1;
logic                             fork2_14_data_out_1_valid;
logic                             fork2_14_data_out_1_ready;
// --------------------------
//   stream_blocks_7_linear1 signals
// --------------------------
logic [stream_blocks_7_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_7_linear1_mdata_in_0        [stream_blocks_7_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_7_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_7_linear1_edata_in_0;
logic                             stream_blocks_7_linear1_data_in_0_valid;
logic                             stream_blocks_7_linear1_data_in_0_ready;
logic [stream_blocks_7_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_7_linear1_mweight        [stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_7_linear1_eweight;
logic                             stream_blocks_7_linear1_weight_valid;
logic                             stream_blocks_7_linear1_weight_ready;
logic [stream_blocks_7_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_7_linear1_mbias        [stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_7_linear1_ebias;
logic                             stream_blocks_7_linear1_bias_valid;
logic                             stream_blocks_7_linear1_bias_ready;
logic [stream_blocks_7_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_7_linear1_mdata_out_0        [stream_blocks_7_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_7_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_7_linear1_edata_out_0;
logic                             stream_blocks_7_linear1_data_out_0_valid;
logic                             stream_blocks_7_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_7_act signals
// --------------------------
logic [stream_blocks_7_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_7_act_mdata_in_0        [stream_blocks_7_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_7_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_7_act_edata_in_0;
logic                             stream_blocks_7_act_data_in_0_valid;
logic                             stream_blocks_7_act_data_in_0_ready;
logic [stream_blocks_7_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_7_act_mdata_out_0        [stream_blocks_7_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_7_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_7_act_edata_out_0;
logic                             stream_blocks_7_act_data_out_0_valid;
logic                             stream_blocks_7_act_data_out_0_ready;
// --------------------------
//   stream_blocks_7_linear2 signals
// --------------------------
logic [stream_blocks_7_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_7_linear2_mdata_in_0        [stream_blocks_7_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_7_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_7_linear2_edata_in_0;
logic                             stream_blocks_7_linear2_data_in_0_valid;
logic                             stream_blocks_7_linear2_data_in_0_ready;
logic [stream_blocks_7_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_7_linear2_mweight        [stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_7_linear2_eweight;
logic                             stream_blocks_7_linear2_weight_valid;
logic                             stream_blocks_7_linear2_weight_ready;
logic [stream_blocks_7_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_7_linear2_mbias        [stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_7_linear2_ebias;
logic                             stream_blocks_7_linear2_bias_valid;
logic                             stream_blocks_7_linear2_bias_ready;
logic [stream_blocks_7_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_7_linear2_mdata_out_0        [stream_blocks_7_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_7_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_7_linear2_edata_out_0;
logic                             stream_blocks_7_linear2_data_out_0_valid;
logic                             stream_blocks_7_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_7_norm1 signals
// --------------------------
logic [stream_blocks_7_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_7_norm1_mdata_in_0        [stream_blocks_7_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_7_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_7_norm1_edata_in_0;
logic                             stream_blocks_7_norm1_data_in_0_valid;
logic                             stream_blocks_7_norm1_data_in_0_ready;
logic [stream_blocks_7_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_7_norm1_mweight        [stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_7_norm1_eweight;
logic                             stream_blocks_7_norm1_weight_valid;
logic                             stream_blocks_7_norm1_weight_ready;
logic [stream_blocks_7_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_7_norm1_mbias        [stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_7_norm1_ebias;
logic                             stream_blocks_7_norm1_bias_valid;
logic                             stream_blocks_7_norm1_bias_ready;
logic [stream_blocks_7_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_7_norm1_mdata_out_0        [stream_blocks_7_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_7_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_7_norm1_edata_out_0;
logic                             stream_blocks_7_norm1_data_out_0_valid;
logic                             stream_blocks_7_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_7_add signals
// --------------------------
logic [stream_blocks_7_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_7_add_mdata_in_0        [stream_blocks_7_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_7_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_7_add_edata_in_0;
logic                             stream_blocks_7_add_data_in_0_valid;
logic                             stream_blocks_7_add_data_in_0_ready;
logic [stream_blocks_7_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_7_add_mdata_in_1        [stream_blocks_7_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_7_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_7_add_edata_in_1;
logic                             stream_blocks_7_add_data_in_1_valid;
logic                             stream_blocks_7_add_data_in_1_ready;
logic [stream_blocks_7_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_7_add_mdata_out_0        [stream_blocks_7_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_7_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_7_add_edata_out_0;
logic                             stream_blocks_7_add_data_out_0_valid;
logic                             stream_blocks_7_add_data_out_0_ready;
// --------------------------
//   fork2_15 signals
// --------------------------
logic [fork2_15_DATA_IN_0_PRECISION_0-1:0]  fork2_15_mdata_in_0        [fork2_15_DATA_IN_0_PARALLELISM_DIM_0*fork2_15_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_15_DATA_IN_0_PRECISION_1-1:0]  fork2_15_edata_in_0;
logic                             fork2_15_data_in_0_valid;
logic                             fork2_15_data_in_0_ready;
logic [fork2_15_DATA_OUT_0_PRECISION_0-1:0]  fork2_15_mdata_out_0        [fork2_15_DATA_OUT_0_PARALLELISM_DIM_0*fork2_15_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_15_DATA_OUT_0_PRECISION_1-1:0]  fork2_15_edata_out_0;
logic                             fork2_15_data_out_0_valid;
logic                             fork2_15_data_out_0_ready;
logic [fork2_15_DATA_OUT_1_PRECISION_0-1:0]  fork2_15_mdata_out_1        [fork2_15_DATA_OUT_1_PARALLELISM_DIM_0*fork2_15_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_15_DATA_OUT_1_PRECISION_1-1:0]  fork2_15_edata_out_1;
logic                             fork2_15_data_out_1_valid;
logic                             fork2_15_data_out_1_ready;
// --------------------------
//   stream_blocks_7_attention signals
// --------------------------
logic [stream_blocks_7_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_7_attention_mdata_in_0        [stream_blocks_7_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_7_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_7_attention_edata_in_0;
logic                             stream_blocks_7_attention_data_in_0_valid;
logic                             stream_blocks_7_attention_data_in_0_ready;
logic [stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_7_attention_mquery_weight        [stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_7_attention_equery_weight;
logic                             stream_blocks_7_attention_query_weight_valid;
logic                             stream_blocks_7_attention_query_weight_ready;
logic [stream_blocks_7_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_7_attention_mquery_bias        [stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_7_attention_equery_bias;
logic                             stream_blocks_7_attention_query_bias_valid;
logic                             stream_blocks_7_attention_query_bias_ready;
logic [stream_blocks_7_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_7_attention_mkey_weight        [stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_7_attention_ekey_weight;
logic                             stream_blocks_7_attention_key_weight_valid;
logic                             stream_blocks_7_attention_key_weight_ready;
logic [stream_blocks_7_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_7_attention_mkey_bias        [stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_7_attention_ekey_bias;
logic                             stream_blocks_7_attention_key_bias_valid;
logic                             stream_blocks_7_attention_key_bias_ready;
logic [stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_7_attention_mvalue_weight        [stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_7_attention_evalue_weight;
logic                             stream_blocks_7_attention_value_weight_valid;
logic                             stream_blocks_7_attention_value_weight_ready;
logic [stream_blocks_7_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_7_attention_mvalue_bias        [stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_7_attention_evalue_bias;
logic                             stream_blocks_7_attention_value_bias_valid;
logic                             stream_blocks_7_attention_value_bias_ready;
logic [stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_7_attention_mproj_weight        [stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_7_attention_eproj_weight;
logic                             stream_blocks_7_attention_proj_weight_valid;
logic                             stream_blocks_7_attention_proj_weight_ready;
logic [stream_blocks_7_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_7_attention_mproj_bias        [stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_7_attention_eproj_bias;
logic                             stream_blocks_7_attention_proj_bias_valid;
logic                             stream_blocks_7_attention_proj_bias_ready;
logic [stream_blocks_7_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_7_attention_mdata_out_0        [stream_blocks_7_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_7_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_7_attention_edata_out_0;
logic                             stream_blocks_7_attention_data_out_0_valid;
logic                             stream_blocks_7_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_7_norm2 signals
// --------------------------
logic [stream_blocks_7_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_7_norm2_mdata_in_0        [stream_blocks_7_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_7_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_7_norm2_edata_in_0;
logic                             stream_blocks_7_norm2_data_in_0_valid;
logic                             stream_blocks_7_norm2_data_in_0_ready;
logic [stream_blocks_7_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_7_norm2_mweight        [stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_7_norm2_eweight;
logic                             stream_blocks_7_norm2_weight_valid;
logic                             stream_blocks_7_norm2_weight_ready;
logic [stream_blocks_7_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_7_norm2_mbias        [stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_7_norm2_ebias;
logic                             stream_blocks_7_norm2_bias_valid;
logic                             stream_blocks_7_norm2_bias_ready;
logic [stream_blocks_7_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_7_norm2_mdata_out_0        [stream_blocks_7_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_7_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_7_norm2_edata_out_0;
logic                             stream_blocks_7_norm2_data_out_0_valid;
logic                             stream_blocks_7_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_7_add_1 signals
// --------------------------
logic [stream_blocks_7_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_7_add_1_mdata_in_0        [stream_blocks_7_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_7_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_7_add_1_edata_in_0;
logic                             stream_blocks_7_add_1_data_in_0_valid;
logic                             stream_blocks_7_add_1_data_in_0_ready;
logic [stream_blocks_7_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_7_add_1_mdata_in_1        [stream_blocks_7_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_7_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_7_add_1_edata_in_1;
logic                             stream_blocks_7_add_1_data_in_1_valid;
logic                             stream_blocks_7_add_1_data_in_1_ready;
logic [stream_blocks_7_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_7_add_1_mdata_out_0        [stream_blocks_7_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_7_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_7_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_7_add_1_edata_out_0;
logic                             stream_blocks_7_add_1_data_out_0_valid;
logic                             stream_blocks_7_add_1_data_out_0_ready;
// --------------------------
//   fork2_16 signals
// --------------------------
logic [fork2_16_DATA_IN_0_PRECISION_0-1:0]  fork2_16_mdata_in_0        [fork2_16_DATA_IN_0_PARALLELISM_DIM_0*fork2_16_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_16_DATA_IN_0_PRECISION_1-1:0]  fork2_16_edata_in_0;
logic                             fork2_16_data_in_0_valid;
logic                             fork2_16_data_in_0_ready;
logic [fork2_16_DATA_OUT_0_PRECISION_0-1:0]  fork2_16_mdata_out_0        [fork2_16_DATA_OUT_0_PARALLELISM_DIM_0*fork2_16_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_16_DATA_OUT_0_PRECISION_1-1:0]  fork2_16_edata_out_0;
logic                             fork2_16_data_out_0_valid;
logic                             fork2_16_data_out_0_ready;
logic [fork2_16_DATA_OUT_1_PRECISION_0-1:0]  fork2_16_mdata_out_1        [fork2_16_DATA_OUT_1_PARALLELISM_DIM_0*fork2_16_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_16_DATA_OUT_1_PRECISION_1-1:0]  fork2_16_edata_out_1;
logic                             fork2_16_data_out_1_valid;
logic                             fork2_16_data_out_1_ready;
// --------------------------
//   stream_blocks_8_linear1 signals
// --------------------------
logic [stream_blocks_8_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_8_linear1_mdata_in_0        [stream_blocks_8_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_8_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_8_linear1_edata_in_0;
logic                             stream_blocks_8_linear1_data_in_0_valid;
logic                             stream_blocks_8_linear1_data_in_0_ready;
logic [stream_blocks_8_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_8_linear1_mweight        [stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_8_linear1_eweight;
logic                             stream_blocks_8_linear1_weight_valid;
logic                             stream_blocks_8_linear1_weight_ready;
logic [stream_blocks_8_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_8_linear1_mbias        [stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_8_linear1_ebias;
logic                             stream_blocks_8_linear1_bias_valid;
logic                             stream_blocks_8_linear1_bias_ready;
logic [stream_blocks_8_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_8_linear1_mdata_out_0        [stream_blocks_8_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_8_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_8_linear1_edata_out_0;
logic                             stream_blocks_8_linear1_data_out_0_valid;
logic                             stream_blocks_8_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_8_act signals
// --------------------------
logic [stream_blocks_8_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_8_act_mdata_in_0        [stream_blocks_8_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_8_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_8_act_edata_in_0;
logic                             stream_blocks_8_act_data_in_0_valid;
logic                             stream_blocks_8_act_data_in_0_ready;
logic [stream_blocks_8_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_8_act_mdata_out_0        [stream_blocks_8_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_8_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_8_act_edata_out_0;
logic                             stream_blocks_8_act_data_out_0_valid;
logic                             stream_blocks_8_act_data_out_0_ready;
// --------------------------
//   stream_blocks_8_linear2 signals
// --------------------------
logic [stream_blocks_8_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_8_linear2_mdata_in_0        [stream_blocks_8_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_8_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_8_linear2_edata_in_0;
logic                             stream_blocks_8_linear2_data_in_0_valid;
logic                             stream_blocks_8_linear2_data_in_0_ready;
logic [stream_blocks_8_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_8_linear2_mweight        [stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_8_linear2_eweight;
logic                             stream_blocks_8_linear2_weight_valid;
logic                             stream_blocks_8_linear2_weight_ready;
logic [stream_blocks_8_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_8_linear2_mbias        [stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_8_linear2_ebias;
logic                             stream_blocks_8_linear2_bias_valid;
logic                             stream_blocks_8_linear2_bias_ready;
logic [stream_blocks_8_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_8_linear2_mdata_out_0        [stream_blocks_8_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_8_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_8_linear2_edata_out_0;
logic                             stream_blocks_8_linear2_data_out_0_valid;
logic                             stream_blocks_8_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_8_norm1 signals
// --------------------------
logic [stream_blocks_8_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_8_norm1_mdata_in_0        [stream_blocks_8_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_8_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_8_norm1_edata_in_0;
logic                             stream_blocks_8_norm1_data_in_0_valid;
logic                             stream_blocks_8_norm1_data_in_0_ready;
logic [stream_blocks_8_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_8_norm1_mweight        [stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_8_norm1_eweight;
logic                             stream_blocks_8_norm1_weight_valid;
logic                             stream_blocks_8_norm1_weight_ready;
logic [stream_blocks_8_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_8_norm1_mbias        [stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_8_norm1_ebias;
logic                             stream_blocks_8_norm1_bias_valid;
logic                             stream_blocks_8_norm1_bias_ready;
logic [stream_blocks_8_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_8_norm1_mdata_out_0        [stream_blocks_8_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_8_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_8_norm1_edata_out_0;
logic                             stream_blocks_8_norm1_data_out_0_valid;
logic                             stream_blocks_8_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_8_add signals
// --------------------------
logic [stream_blocks_8_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_8_add_mdata_in_0        [stream_blocks_8_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_8_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_8_add_edata_in_0;
logic                             stream_blocks_8_add_data_in_0_valid;
logic                             stream_blocks_8_add_data_in_0_ready;
logic [stream_blocks_8_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_8_add_mdata_in_1        [stream_blocks_8_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_8_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_8_add_edata_in_1;
logic                             stream_blocks_8_add_data_in_1_valid;
logic                             stream_blocks_8_add_data_in_1_ready;
logic [stream_blocks_8_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_8_add_mdata_out_0        [stream_blocks_8_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_8_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_8_add_edata_out_0;
logic                             stream_blocks_8_add_data_out_0_valid;
logic                             stream_blocks_8_add_data_out_0_ready;
// --------------------------
//   fork2_17 signals
// --------------------------
logic [fork2_17_DATA_IN_0_PRECISION_0-1:0]  fork2_17_mdata_in_0        [fork2_17_DATA_IN_0_PARALLELISM_DIM_0*fork2_17_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_17_DATA_IN_0_PRECISION_1-1:0]  fork2_17_edata_in_0;
logic                             fork2_17_data_in_0_valid;
logic                             fork2_17_data_in_0_ready;
logic [fork2_17_DATA_OUT_0_PRECISION_0-1:0]  fork2_17_mdata_out_0        [fork2_17_DATA_OUT_0_PARALLELISM_DIM_0*fork2_17_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_17_DATA_OUT_0_PRECISION_1-1:0]  fork2_17_edata_out_0;
logic                             fork2_17_data_out_0_valid;
logic                             fork2_17_data_out_0_ready;
logic [fork2_17_DATA_OUT_1_PRECISION_0-1:0]  fork2_17_mdata_out_1        [fork2_17_DATA_OUT_1_PARALLELISM_DIM_0*fork2_17_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_17_DATA_OUT_1_PRECISION_1-1:0]  fork2_17_edata_out_1;
logic                             fork2_17_data_out_1_valid;
logic                             fork2_17_data_out_1_ready;
// --------------------------
//   stream_blocks_8_attention signals
// --------------------------
logic [stream_blocks_8_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_8_attention_mdata_in_0        [stream_blocks_8_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_8_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_8_attention_edata_in_0;
logic                             stream_blocks_8_attention_data_in_0_valid;
logic                             stream_blocks_8_attention_data_in_0_ready;
logic [stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_8_attention_mquery_weight        [stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_8_attention_equery_weight;
logic                             stream_blocks_8_attention_query_weight_valid;
logic                             stream_blocks_8_attention_query_weight_ready;
logic [stream_blocks_8_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_8_attention_mquery_bias        [stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_8_attention_equery_bias;
logic                             stream_blocks_8_attention_query_bias_valid;
logic                             stream_blocks_8_attention_query_bias_ready;
logic [stream_blocks_8_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_8_attention_mkey_weight        [stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_8_attention_ekey_weight;
logic                             stream_blocks_8_attention_key_weight_valid;
logic                             stream_blocks_8_attention_key_weight_ready;
logic [stream_blocks_8_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_8_attention_mkey_bias        [stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_8_attention_ekey_bias;
logic                             stream_blocks_8_attention_key_bias_valid;
logic                             stream_blocks_8_attention_key_bias_ready;
logic [stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_8_attention_mvalue_weight        [stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_8_attention_evalue_weight;
logic                             stream_blocks_8_attention_value_weight_valid;
logic                             stream_blocks_8_attention_value_weight_ready;
logic [stream_blocks_8_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_8_attention_mvalue_bias        [stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_8_attention_evalue_bias;
logic                             stream_blocks_8_attention_value_bias_valid;
logic                             stream_blocks_8_attention_value_bias_ready;
logic [stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_8_attention_mproj_weight        [stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_8_attention_eproj_weight;
logic                             stream_blocks_8_attention_proj_weight_valid;
logic                             stream_blocks_8_attention_proj_weight_ready;
logic [stream_blocks_8_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_8_attention_mproj_bias        [stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_8_attention_eproj_bias;
logic                             stream_blocks_8_attention_proj_bias_valid;
logic                             stream_blocks_8_attention_proj_bias_ready;
logic [stream_blocks_8_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_8_attention_mdata_out_0        [stream_blocks_8_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_8_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_8_attention_edata_out_0;
logic                             stream_blocks_8_attention_data_out_0_valid;
logic                             stream_blocks_8_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_8_norm2 signals
// --------------------------
logic [stream_blocks_8_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_8_norm2_mdata_in_0        [stream_blocks_8_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_8_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_8_norm2_edata_in_0;
logic                             stream_blocks_8_norm2_data_in_0_valid;
logic                             stream_blocks_8_norm2_data_in_0_ready;
logic [stream_blocks_8_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_8_norm2_mweight        [stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_8_norm2_eweight;
logic                             stream_blocks_8_norm2_weight_valid;
logic                             stream_blocks_8_norm2_weight_ready;
logic [stream_blocks_8_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_8_norm2_mbias        [stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_8_norm2_ebias;
logic                             stream_blocks_8_norm2_bias_valid;
logic                             stream_blocks_8_norm2_bias_ready;
logic [stream_blocks_8_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_8_norm2_mdata_out_0        [stream_blocks_8_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_8_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_8_norm2_edata_out_0;
logic                             stream_blocks_8_norm2_data_out_0_valid;
logic                             stream_blocks_8_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_8_add_1 signals
// --------------------------
logic [stream_blocks_8_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_8_add_1_mdata_in_0        [stream_blocks_8_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_8_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_8_add_1_edata_in_0;
logic                             stream_blocks_8_add_1_data_in_0_valid;
logic                             stream_blocks_8_add_1_data_in_0_ready;
logic [stream_blocks_8_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_8_add_1_mdata_in_1        [stream_blocks_8_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_8_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_8_add_1_edata_in_1;
logic                             stream_blocks_8_add_1_data_in_1_valid;
logic                             stream_blocks_8_add_1_data_in_1_ready;
logic [stream_blocks_8_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_8_add_1_mdata_out_0        [stream_blocks_8_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_8_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_8_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_8_add_1_edata_out_0;
logic                             stream_blocks_8_add_1_data_out_0_valid;
logic                             stream_blocks_8_add_1_data_out_0_ready;
// --------------------------
//   fork2_18 signals
// --------------------------
logic [fork2_18_DATA_IN_0_PRECISION_0-1:0]  fork2_18_mdata_in_0        [fork2_18_DATA_IN_0_PARALLELISM_DIM_0*fork2_18_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_18_DATA_IN_0_PRECISION_1-1:0]  fork2_18_edata_in_0;
logic                             fork2_18_data_in_0_valid;
logic                             fork2_18_data_in_0_ready;
logic [fork2_18_DATA_OUT_0_PRECISION_0-1:0]  fork2_18_mdata_out_0        [fork2_18_DATA_OUT_0_PARALLELISM_DIM_0*fork2_18_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_18_DATA_OUT_0_PRECISION_1-1:0]  fork2_18_edata_out_0;
logic                             fork2_18_data_out_0_valid;
logic                             fork2_18_data_out_0_ready;
logic [fork2_18_DATA_OUT_1_PRECISION_0-1:0]  fork2_18_mdata_out_1        [fork2_18_DATA_OUT_1_PARALLELISM_DIM_0*fork2_18_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_18_DATA_OUT_1_PRECISION_1-1:0]  fork2_18_edata_out_1;
logic                             fork2_18_data_out_1_valid;
logic                             fork2_18_data_out_1_ready;
// --------------------------
//   stream_blocks_9_linear1 signals
// --------------------------
logic [stream_blocks_9_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_9_linear1_mdata_in_0        [stream_blocks_9_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_9_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_9_linear1_edata_in_0;
logic                             stream_blocks_9_linear1_data_in_0_valid;
logic                             stream_blocks_9_linear1_data_in_0_ready;
logic [stream_blocks_9_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_9_linear1_mweight        [stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_9_linear1_eweight;
logic                             stream_blocks_9_linear1_weight_valid;
logic                             stream_blocks_9_linear1_weight_ready;
logic [stream_blocks_9_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_9_linear1_mbias        [stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_9_linear1_ebias;
logic                             stream_blocks_9_linear1_bias_valid;
logic                             stream_blocks_9_linear1_bias_ready;
logic [stream_blocks_9_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_9_linear1_mdata_out_0        [stream_blocks_9_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_9_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_9_linear1_edata_out_0;
logic                             stream_blocks_9_linear1_data_out_0_valid;
logic                             stream_blocks_9_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_9_act signals
// --------------------------
logic [stream_blocks_9_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_9_act_mdata_in_0        [stream_blocks_9_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_9_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_9_act_edata_in_0;
logic                             stream_blocks_9_act_data_in_0_valid;
logic                             stream_blocks_9_act_data_in_0_ready;
logic [stream_blocks_9_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_9_act_mdata_out_0        [stream_blocks_9_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_9_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_9_act_edata_out_0;
logic                             stream_blocks_9_act_data_out_0_valid;
logic                             stream_blocks_9_act_data_out_0_ready;
// --------------------------
//   stream_blocks_9_linear2 signals
// --------------------------
logic [stream_blocks_9_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_9_linear2_mdata_in_0        [stream_blocks_9_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_9_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_9_linear2_edata_in_0;
logic                             stream_blocks_9_linear2_data_in_0_valid;
logic                             stream_blocks_9_linear2_data_in_0_ready;
logic [stream_blocks_9_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_9_linear2_mweight        [stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_9_linear2_eweight;
logic                             stream_blocks_9_linear2_weight_valid;
logic                             stream_blocks_9_linear2_weight_ready;
logic [stream_blocks_9_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_9_linear2_mbias        [stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_9_linear2_ebias;
logic                             stream_blocks_9_linear2_bias_valid;
logic                             stream_blocks_9_linear2_bias_ready;
logic [stream_blocks_9_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_9_linear2_mdata_out_0        [stream_blocks_9_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_9_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_9_linear2_edata_out_0;
logic                             stream_blocks_9_linear2_data_out_0_valid;
logic                             stream_blocks_9_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_9_norm1 signals
// --------------------------
logic [stream_blocks_9_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_9_norm1_mdata_in_0        [stream_blocks_9_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_9_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_9_norm1_edata_in_0;
logic                             stream_blocks_9_norm1_data_in_0_valid;
logic                             stream_blocks_9_norm1_data_in_0_ready;
logic [stream_blocks_9_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_9_norm1_mweight        [stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_9_norm1_eweight;
logic                             stream_blocks_9_norm1_weight_valid;
logic                             stream_blocks_9_norm1_weight_ready;
logic [stream_blocks_9_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_9_norm1_mbias        [stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_9_norm1_ebias;
logic                             stream_blocks_9_norm1_bias_valid;
logic                             stream_blocks_9_norm1_bias_ready;
logic [stream_blocks_9_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_9_norm1_mdata_out_0        [stream_blocks_9_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_9_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_9_norm1_edata_out_0;
logic                             stream_blocks_9_norm1_data_out_0_valid;
logic                             stream_blocks_9_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_9_add signals
// --------------------------
logic [stream_blocks_9_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_9_add_mdata_in_0        [stream_blocks_9_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_9_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_9_add_edata_in_0;
logic                             stream_blocks_9_add_data_in_0_valid;
logic                             stream_blocks_9_add_data_in_0_ready;
logic [stream_blocks_9_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_9_add_mdata_in_1        [stream_blocks_9_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_9_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_9_add_edata_in_1;
logic                             stream_blocks_9_add_data_in_1_valid;
logic                             stream_blocks_9_add_data_in_1_ready;
logic [stream_blocks_9_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_9_add_mdata_out_0        [stream_blocks_9_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_9_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_9_add_edata_out_0;
logic                             stream_blocks_9_add_data_out_0_valid;
logic                             stream_blocks_9_add_data_out_0_ready;
// --------------------------
//   fork2_19 signals
// --------------------------
logic [fork2_19_DATA_IN_0_PRECISION_0-1:0]  fork2_19_mdata_in_0        [fork2_19_DATA_IN_0_PARALLELISM_DIM_0*fork2_19_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_19_DATA_IN_0_PRECISION_1-1:0]  fork2_19_edata_in_0;
logic                             fork2_19_data_in_0_valid;
logic                             fork2_19_data_in_0_ready;
logic [fork2_19_DATA_OUT_0_PRECISION_0-1:0]  fork2_19_mdata_out_0        [fork2_19_DATA_OUT_0_PARALLELISM_DIM_0*fork2_19_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_19_DATA_OUT_0_PRECISION_1-1:0]  fork2_19_edata_out_0;
logic                             fork2_19_data_out_0_valid;
logic                             fork2_19_data_out_0_ready;
logic [fork2_19_DATA_OUT_1_PRECISION_0-1:0]  fork2_19_mdata_out_1        [fork2_19_DATA_OUT_1_PARALLELISM_DIM_0*fork2_19_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_19_DATA_OUT_1_PRECISION_1-1:0]  fork2_19_edata_out_1;
logic                             fork2_19_data_out_1_valid;
logic                             fork2_19_data_out_1_ready;
// --------------------------
//   stream_blocks_9_attention signals
// --------------------------
logic [stream_blocks_9_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_9_attention_mdata_in_0        [stream_blocks_9_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_9_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_9_attention_edata_in_0;
logic                             stream_blocks_9_attention_data_in_0_valid;
logic                             stream_blocks_9_attention_data_in_0_ready;
logic [stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_9_attention_mquery_weight        [stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_9_attention_equery_weight;
logic                             stream_blocks_9_attention_query_weight_valid;
logic                             stream_blocks_9_attention_query_weight_ready;
logic [stream_blocks_9_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_9_attention_mquery_bias        [stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_9_attention_equery_bias;
logic                             stream_blocks_9_attention_query_bias_valid;
logic                             stream_blocks_9_attention_query_bias_ready;
logic [stream_blocks_9_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_9_attention_mkey_weight        [stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_9_attention_ekey_weight;
logic                             stream_blocks_9_attention_key_weight_valid;
logic                             stream_blocks_9_attention_key_weight_ready;
logic [stream_blocks_9_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_9_attention_mkey_bias        [stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_9_attention_ekey_bias;
logic                             stream_blocks_9_attention_key_bias_valid;
logic                             stream_blocks_9_attention_key_bias_ready;
logic [stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_9_attention_mvalue_weight        [stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_9_attention_evalue_weight;
logic                             stream_blocks_9_attention_value_weight_valid;
logic                             stream_blocks_9_attention_value_weight_ready;
logic [stream_blocks_9_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_9_attention_mvalue_bias        [stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_9_attention_evalue_bias;
logic                             stream_blocks_9_attention_value_bias_valid;
logic                             stream_blocks_9_attention_value_bias_ready;
logic [stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_9_attention_mproj_weight        [stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_9_attention_eproj_weight;
logic                             stream_blocks_9_attention_proj_weight_valid;
logic                             stream_blocks_9_attention_proj_weight_ready;
logic [stream_blocks_9_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_9_attention_mproj_bias        [stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_9_attention_eproj_bias;
logic                             stream_blocks_9_attention_proj_bias_valid;
logic                             stream_blocks_9_attention_proj_bias_ready;
logic [stream_blocks_9_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_9_attention_mdata_out_0        [stream_blocks_9_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_9_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_9_attention_edata_out_0;
logic                             stream_blocks_9_attention_data_out_0_valid;
logic                             stream_blocks_9_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_9_norm2 signals
// --------------------------
logic [stream_blocks_9_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_9_norm2_mdata_in_0        [stream_blocks_9_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_9_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_9_norm2_edata_in_0;
logic                             stream_blocks_9_norm2_data_in_0_valid;
logic                             stream_blocks_9_norm2_data_in_0_ready;
logic [stream_blocks_9_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_9_norm2_mweight        [stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_9_norm2_eweight;
logic                             stream_blocks_9_norm2_weight_valid;
logic                             stream_blocks_9_norm2_weight_ready;
logic [stream_blocks_9_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_9_norm2_mbias        [stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_9_norm2_ebias;
logic                             stream_blocks_9_norm2_bias_valid;
logic                             stream_blocks_9_norm2_bias_ready;
logic [stream_blocks_9_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_9_norm2_mdata_out_0        [stream_blocks_9_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_9_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_9_norm2_edata_out_0;
logic                             stream_blocks_9_norm2_data_out_0_valid;
logic                             stream_blocks_9_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_9_add_1 signals
// --------------------------
logic [stream_blocks_9_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_9_add_1_mdata_in_0        [stream_blocks_9_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_9_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_9_add_1_edata_in_0;
logic                             stream_blocks_9_add_1_data_in_0_valid;
logic                             stream_blocks_9_add_1_data_in_0_ready;
logic [stream_blocks_9_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_9_add_1_mdata_in_1        [stream_blocks_9_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_9_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_9_add_1_edata_in_1;
logic                             stream_blocks_9_add_1_data_in_1_valid;
logic                             stream_blocks_9_add_1_data_in_1_ready;
logic [stream_blocks_9_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_9_add_1_mdata_out_0        [stream_blocks_9_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_9_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_9_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_9_add_1_edata_out_0;
logic                             stream_blocks_9_add_1_data_out_0_valid;
logic                             stream_blocks_9_add_1_data_out_0_ready;
// --------------------------
//   fork2_20 signals
// --------------------------
logic [fork2_20_DATA_IN_0_PRECISION_0-1:0]  fork2_20_mdata_in_0        [fork2_20_DATA_IN_0_PARALLELISM_DIM_0*fork2_20_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_20_DATA_IN_0_PRECISION_1-1:0]  fork2_20_edata_in_0;
logic                             fork2_20_data_in_0_valid;
logic                             fork2_20_data_in_0_ready;
logic [fork2_20_DATA_OUT_0_PRECISION_0-1:0]  fork2_20_mdata_out_0        [fork2_20_DATA_OUT_0_PARALLELISM_DIM_0*fork2_20_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_20_DATA_OUT_0_PRECISION_1-1:0]  fork2_20_edata_out_0;
logic                             fork2_20_data_out_0_valid;
logic                             fork2_20_data_out_0_ready;
logic [fork2_20_DATA_OUT_1_PRECISION_0-1:0]  fork2_20_mdata_out_1        [fork2_20_DATA_OUT_1_PARALLELISM_DIM_0*fork2_20_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_20_DATA_OUT_1_PRECISION_1-1:0]  fork2_20_edata_out_1;
logic                             fork2_20_data_out_1_valid;
logic                             fork2_20_data_out_1_ready;
// --------------------------
//   stream_blocks_10_linear1 signals
// --------------------------
logic [stream_blocks_10_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_10_linear1_mdata_in_0        [stream_blocks_10_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_10_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_10_linear1_edata_in_0;
logic                             stream_blocks_10_linear1_data_in_0_valid;
logic                             stream_blocks_10_linear1_data_in_0_ready;
logic [stream_blocks_10_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_10_linear1_mweight        [stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_10_linear1_eweight;
logic                             stream_blocks_10_linear1_weight_valid;
logic                             stream_blocks_10_linear1_weight_ready;
logic [stream_blocks_10_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_10_linear1_mbias        [stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_10_linear1_ebias;
logic                             stream_blocks_10_linear1_bias_valid;
logic                             stream_blocks_10_linear1_bias_ready;
logic [stream_blocks_10_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_10_linear1_mdata_out_0        [stream_blocks_10_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_10_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_10_linear1_edata_out_0;
logic                             stream_blocks_10_linear1_data_out_0_valid;
logic                             stream_blocks_10_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_10_act signals
// --------------------------
logic [stream_blocks_10_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_10_act_mdata_in_0        [stream_blocks_10_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_10_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_10_act_edata_in_0;
logic                             stream_blocks_10_act_data_in_0_valid;
logic                             stream_blocks_10_act_data_in_0_ready;
logic [stream_blocks_10_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_10_act_mdata_out_0        [stream_blocks_10_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_10_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_10_act_edata_out_0;
logic                             stream_blocks_10_act_data_out_0_valid;
logic                             stream_blocks_10_act_data_out_0_ready;
// --------------------------
//   stream_blocks_10_linear2 signals
// --------------------------
logic [stream_blocks_10_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_10_linear2_mdata_in_0        [stream_blocks_10_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_10_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_10_linear2_edata_in_0;
logic                             stream_blocks_10_linear2_data_in_0_valid;
logic                             stream_blocks_10_linear2_data_in_0_ready;
logic [stream_blocks_10_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_10_linear2_mweight        [stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_10_linear2_eweight;
logic                             stream_blocks_10_linear2_weight_valid;
logic                             stream_blocks_10_linear2_weight_ready;
logic [stream_blocks_10_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_10_linear2_mbias        [stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_10_linear2_ebias;
logic                             stream_blocks_10_linear2_bias_valid;
logic                             stream_blocks_10_linear2_bias_ready;
logic [stream_blocks_10_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_10_linear2_mdata_out_0        [stream_blocks_10_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_10_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_10_linear2_edata_out_0;
logic                             stream_blocks_10_linear2_data_out_0_valid;
logic                             stream_blocks_10_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_10_norm1 signals
// --------------------------
logic [stream_blocks_10_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_10_norm1_mdata_in_0        [stream_blocks_10_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_10_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_10_norm1_edata_in_0;
logic                             stream_blocks_10_norm1_data_in_0_valid;
logic                             stream_blocks_10_norm1_data_in_0_ready;
logic [stream_blocks_10_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_10_norm1_mweight        [stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_10_norm1_eweight;
logic                             stream_blocks_10_norm1_weight_valid;
logic                             stream_blocks_10_norm1_weight_ready;
logic [stream_blocks_10_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_10_norm1_mbias        [stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_10_norm1_ebias;
logic                             stream_blocks_10_norm1_bias_valid;
logic                             stream_blocks_10_norm1_bias_ready;
logic [stream_blocks_10_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_10_norm1_mdata_out_0        [stream_blocks_10_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_10_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_10_norm1_edata_out_0;
logic                             stream_blocks_10_norm1_data_out_0_valid;
logic                             stream_blocks_10_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_10_add signals
// --------------------------
logic [stream_blocks_10_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_10_add_mdata_in_0        [stream_blocks_10_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_10_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_10_add_edata_in_0;
logic                             stream_blocks_10_add_data_in_0_valid;
logic                             stream_blocks_10_add_data_in_0_ready;
logic [stream_blocks_10_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_10_add_mdata_in_1        [stream_blocks_10_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_10_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_10_add_edata_in_1;
logic                             stream_blocks_10_add_data_in_1_valid;
logic                             stream_blocks_10_add_data_in_1_ready;
logic [stream_blocks_10_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_10_add_mdata_out_0        [stream_blocks_10_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_10_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_10_add_edata_out_0;
logic                             stream_blocks_10_add_data_out_0_valid;
logic                             stream_blocks_10_add_data_out_0_ready;
// --------------------------
//   fork2_21 signals
// --------------------------
logic [fork2_21_DATA_IN_0_PRECISION_0-1:0]  fork2_21_mdata_in_0        [fork2_21_DATA_IN_0_PARALLELISM_DIM_0*fork2_21_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_21_DATA_IN_0_PRECISION_1-1:0]  fork2_21_edata_in_0;
logic                             fork2_21_data_in_0_valid;
logic                             fork2_21_data_in_0_ready;
logic [fork2_21_DATA_OUT_0_PRECISION_0-1:0]  fork2_21_mdata_out_0        [fork2_21_DATA_OUT_0_PARALLELISM_DIM_0*fork2_21_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_21_DATA_OUT_0_PRECISION_1-1:0]  fork2_21_edata_out_0;
logic                             fork2_21_data_out_0_valid;
logic                             fork2_21_data_out_0_ready;
logic [fork2_21_DATA_OUT_1_PRECISION_0-1:0]  fork2_21_mdata_out_1        [fork2_21_DATA_OUT_1_PARALLELISM_DIM_0*fork2_21_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_21_DATA_OUT_1_PRECISION_1-1:0]  fork2_21_edata_out_1;
logic                             fork2_21_data_out_1_valid;
logic                             fork2_21_data_out_1_ready;
// --------------------------
//   stream_blocks_10_attention signals
// --------------------------
logic [stream_blocks_10_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_10_attention_mdata_in_0        [stream_blocks_10_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_10_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_10_attention_edata_in_0;
logic                             stream_blocks_10_attention_data_in_0_valid;
logic                             stream_blocks_10_attention_data_in_0_ready;
logic [stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_10_attention_mquery_weight        [stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_10_attention_equery_weight;
logic                             stream_blocks_10_attention_query_weight_valid;
logic                             stream_blocks_10_attention_query_weight_ready;
logic [stream_blocks_10_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_10_attention_mquery_bias        [stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_10_attention_equery_bias;
logic                             stream_blocks_10_attention_query_bias_valid;
logic                             stream_blocks_10_attention_query_bias_ready;
logic [stream_blocks_10_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_10_attention_mkey_weight        [stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_10_attention_ekey_weight;
logic                             stream_blocks_10_attention_key_weight_valid;
logic                             stream_blocks_10_attention_key_weight_ready;
logic [stream_blocks_10_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_10_attention_mkey_bias        [stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_10_attention_ekey_bias;
logic                             stream_blocks_10_attention_key_bias_valid;
logic                             stream_blocks_10_attention_key_bias_ready;
logic [stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_10_attention_mvalue_weight        [stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_10_attention_evalue_weight;
logic                             stream_blocks_10_attention_value_weight_valid;
logic                             stream_blocks_10_attention_value_weight_ready;
logic [stream_blocks_10_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_10_attention_mvalue_bias        [stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_10_attention_evalue_bias;
logic                             stream_blocks_10_attention_value_bias_valid;
logic                             stream_blocks_10_attention_value_bias_ready;
logic [stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_10_attention_mproj_weight        [stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_10_attention_eproj_weight;
logic                             stream_blocks_10_attention_proj_weight_valid;
logic                             stream_blocks_10_attention_proj_weight_ready;
logic [stream_blocks_10_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_10_attention_mproj_bias        [stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_10_attention_eproj_bias;
logic                             stream_blocks_10_attention_proj_bias_valid;
logic                             stream_blocks_10_attention_proj_bias_ready;
logic [stream_blocks_10_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_10_attention_mdata_out_0        [stream_blocks_10_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_10_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_10_attention_edata_out_0;
logic                             stream_blocks_10_attention_data_out_0_valid;
logic                             stream_blocks_10_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_10_norm2 signals
// --------------------------
logic [stream_blocks_10_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_10_norm2_mdata_in_0        [stream_blocks_10_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_10_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_10_norm2_edata_in_0;
logic                             stream_blocks_10_norm2_data_in_0_valid;
logic                             stream_blocks_10_norm2_data_in_0_ready;
logic [stream_blocks_10_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_10_norm2_mweight        [stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_10_norm2_eweight;
logic                             stream_blocks_10_norm2_weight_valid;
logic                             stream_blocks_10_norm2_weight_ready;
logic [stream_blocks_10_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_10_norm2_mbias        [stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_10_norm2_ebias;
logic                             stream_blocks_10_norm2_bias_valid;
logic                             stream_blocks_10_norm2_bias_ready;
logic [stream_blocks_10_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_10_norm2_mdata_out_0        [stream_blocks_10_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_10_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_10_norm2_edata_out_0;
logic                             stream_blocks_10_norm2_data_out_0_valid;
logic                             stream_blocks_10_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_10_add_1 signals
// --------------------------
logic [stream_blocks_10_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_10_add_1_mdata_in_0        [stream_blocks_10_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_10_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_10_add_1_edata_in_0;
logic                             stream_blocks_10_add_1_data_in_0_valid;
logic                             stream_blocks_10_add_1_data_in_0_ready;
logic [stream_blocks_10_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_10_add_1_mdata_in_1        [stream_blocks_10_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_10_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_10_add_1_edata_in_1;
logic                             stream_blocks_10_add_1_data_in_1_valid;
logic                             stream_blocks_10_add_1_data_in_1_ready;
logic [stream_blocks_10_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_10_add_1_mdata_out_0        [stream_blocks_10_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_10_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_10_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_10_add_1_edata_out_0;
logic                             stream_blocks_10_add_1_data_out_0_valid;
logic                             stream_blocks_10_add_1_data_out_0_ready;
// --------------------------
//   fork2_22 signals
// --------------------------
logic [fork2_22_DATA_IN_0_PRECISION_0-1:0]  fork2_22_mdata_in_0        [fork2_22_DATA_IN_0_PARALLELISM_DIM_0*fork2_22_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_22_DATA_IN_0_PRECISION_1-1:0]  fork2_22_edata_in_0;
logic                             fork2_22_data_in_0_valid;
logic                             fork2_22_data_in_0_ready;
logic [fork2_22_DATA_OUT_0_PRECISION_0-1:0]  fork2_22_mdata_out_0        [fork2_22_DATA_OUT_0_PARALLELISM_DIM_0*fork2_22_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_22_DATA_OUT_0_PRECISION_1-1:0]  fork2_22_edata_out_0;
logic                             fork2_22_data_out_0_valid;
logic                             fork2_22_data_out_0_ready;
logic [fork2_22_DATA_OUT_1_PRECISION_0-1:0]  fork2_22_mdata_out_1        [fork2_22_DATA_OUT_1_PARALLELISM_DIM_0*fork2_22_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_22_DATA_OUT_1_PRECISION_1-1:0]  fork2_22_edata_out_1;
logic                             fork2_22_data_out_1_valid;
logic                             fork2_22_data_out_1_ready;
// --------------------------
//   stream_blocks_11_linear1 signals
// --------------------------
logic [stream_blocks_11_linear1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_11_linear1_mdata_in_0        [stream_blocks_11_linear1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_11_linear1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_linear1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_11_linear1_edata_in_0;
logic                             stream_blocks_11_linear1_data_in_0_valid;
logic                             stream_blocks_11_linear1_data_in_0_ready;
logic [stream_blocks_11_linear1_WEIGHT_PRECISION_0-1:0]  stream_blocks_11_linear1_mweight        [stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_linear1_WEIGHT_PRECISION_1-1:0]  stream_blocks_11_linear1_eweight;
logic                             stream_blocks_11_linear1_weight_valid;
logic                             stream_blocks_11_linear1_weight_ready;
logic [stream_blocks_11_linear1_BIAS_PRECISION_0-1:0]  stream_blocks_11_linear1_mbias        [stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_0*stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_linear1_BIAS_PRECISION_1-1:0]  stream_blocks_11_linear1_ebias;
logic                             stream_blocks_11_linear1_bias_valid;
logic                             stream_blocks_11_linear1_bias_ready;
logic [stream_blocks_11_linear1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_11_linear1_mdata_out_0        [stream_blocks_11_linear1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_11_linear1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_linear1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_11_linear1_edata_out_0;
logic                             stream_blocks_11_linear1_data_out_0_valid;
logic                             stream_blocks_11_linear1_data_out_0_ready;
// --------------------------
//   stream_blocks_11_act signals
// --------------------------
logic [stream_blocks_11_act_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_11_act_mdata_in_0        [stream_blocks_11_act_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_11_act_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_act_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_11_act_edata_in_0;
logic                             stream_blocks_11_act_data_in_0_valid;
logic                             stream_blocks_11_act_data_in_0_ready;
logic [stream_blocks_11_act_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_11_act_mdata_out_0        [stream_blocks_11_act_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_11_act_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_act_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_11_act_edata_out_0;
logic                             stream_blocks_11_act_data_out_0_valid;
logic                             stream_blocks_11_act_data_out_0_ready;
// --------------------------
//   stream_blocks_11_linear2 signals
// --------------------------
logic [stream_blocks_11_linear2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_11_linear2_mdata_in_0        [stream_blocks_11_linear2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_11_linear2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_linear2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_11_linear2_edata_in_0;
logic                             stream_blocks_11_linear2_data_in_0_valid;
logic                             stream_blocks_11_linear2_data_in_0_ready;
logic [stream_blocks_11_linear2_WEIGHT_PRECISION_0-1:0]  stream_blocks_11_linear2_mweight        [stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_linear2_WEIGHT_PRECISION_1-1:0]  stream_blocks_11_linear2_eweight;
logic                             stream_blocks_11_linear2_weight_valid;
logic                             stream_blocks_11_linear2_weight_ready;
logic [stream_blocks_11_linear2_BIAS_PRECISION_0-1:0]  stream_blocks_11_linear2_mbias        [stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_0*stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_linear2_BIAS_PRECISION_1-1:0]  stream_blocks_11_linear2_ebias;
logic                             stream_blocks_11_linear2_bias_valid;
logic                             stream_blocks_11_linear2_bias_ready;
logic [stream_blocks_11_linear2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_11_linear2_mdata_out_0        [stream_blocks_11_linear2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_11_linear2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_linear2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_11_linear2_edata_out_0;
logic                             stream_blocks_11_linear2_data_out_0_valid;
logic                             stream_blocks_11_linear2_data_out_0_ready;
// --------------------------
//   stream_blocks_11_norm1 signals
// --------------------------
logic [stream_blocks_11_norm1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_11_norm1_mdata_in_0        [stream_blocks_11_norm1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_11_norm1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_norm1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_11_norm1_edata_in_0;
logic                             stream_blocks_11_norm1_data_in_0_valid;
logic                             stream_blocks_11_norm1_data_in_0_ready;
logic [stream_blocks_11_norm1_WEIGHT_PRECISION_0-1:0]  stream_blocks_11_norm1_mweight        [stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_0*stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_norm1_WEIGHT_PRECISION_1-1:0]  stream_blocks_11_norm1_eweight;
logic                             stream_blocks_11_norm1_weight_valid;
logic                             stream_blocks_11_norm1_weight_ready;
logic [stream_blocks_11_norm1_BIAS_PRECISION_0-1:0]  stream_blocks_11_norm1_mbias        [stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_0*stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_norm1_BIAS_PRECISION_1-1:0]  stream_blocks_11_norm1_ebias;
logic                             stream_blocks_11_norm1_bias_valid;
logic                             stream_blocks_11_norm1_bias_ready;
logic [stream_blocks_11_norm1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_11_norm1_mdata_out_0        [stream_blocks_11_norm1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_11_norm1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_norm1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_11_norm1_edata_out_0;
logic                             stream_blocks_11_norm1_data_out_0_valid;
logic                             stream_blocks_11_norm1_data_out_0_ready;
// --------------------------
//   stream_blocks_11_add signals
// --------------------------
logic [stream_blocks_11_add_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_11_add_mdata_in_0        [stream_blocks_11_add_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_11_add_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_add_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_11_add_edata_in_0;
logic                             stream_blocks_11_add_data_in_0_valid;
logic                             stream_blocks_11_add_data_in_0_ready;
logic [stream_blocks_11_add_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_11_add_mdata_in_1        [stream_blocks_11_add_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_11_add_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_add_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_11_add_edata_in_1;
logic                             stream_blocks_11_add_data_in_1_valid;
logic                             stream_blocks_11_add_data_in_1_ready;
logic [stream_blocks_11_add_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_11_add_mdata_out_0        [stream_blocks_11_add_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_11_add_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_add_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_11_add_edata_out_0;
logic                             stream_blocks_11_add_data_out_0_valid;
logic                             stream_blocks_11_add_data_out_0_ready;
// --------------------------
//   fork2_23 signals
// --------------------------
logic [fork2_23_DATA_IN_0_PRECISION_0-1:0]  fork2_23_mdata_in_0        [fork2_23_DATA_IN_0_PARALLELISM_DIM_0*fork2_23_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [fork2_23_DATA_IN_0_PRECISION_1-1:0]  fork2_23_edata_in_0;
logic                             fork2_23_data_in_0_valid;
logic                             fork2_23_data_in_0_ready;
logic [fork2_23_DATA_OUT_0_PRECISION_0-1:0]  fork2_23_mdata_out_0        [fork2_23_DATA_OUT_0_PARALLELISM_DIM_0*fork2_23_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [fork2_23_DATA_OUT_0_PRECISION_1-1:0]  fork2_23_edata_out_0;
logic                             fork2_23_data_out_0_valid;
logic                             fork2_23_data_out_0_ready;
logic [fork2_23_DATA_OUT_1_PRECISION_0-1:0]  fork2_23_mdata_out_1        [fork2_23_DATA_OUT_1_PARALLELISM_DIM_0*fork2_23_DATA_OUT_1_PARALLELISM_DIM_1-1:0];
logic [fork2_23_DATA_OUT_1_PRECISION_1-1:0]  fork2_23_edata_out_1;
logic                             fork2_23_data_out_1_valid;
logic                             fork2_23_data_out_1_ready;
// --------------------------
//   stream_blocks_11_attention signals
// --------------------------
logic [stream_blocks_11_attention_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_11_attention_mdata_in_0        [stream_blocks_11_attention_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_11_attention_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_11_attention_edata_in_0;
logic                             stream_blocks_11_attention_data_in_0_valid;
logic                             stream_blocks_11_attention_data_in_0_ready;
logic [stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_0-1:0]  stream_blocks_11_attention_mquery_weight        [stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_1-1:0]  stream_blocks_11_attention_equery_weight;
logic                             stream_blocks_11_attention_query_weight_valid;
logic                             stream_blocks_11_attention_query_weight_ready;
logic [stream_blocks_11_attention_QUERY_BIAS_PRECISION_0-1:0]  stream_blocks_11_attention_mquery_bias        [stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_0*stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_QUERY_BIAS_PRECISION_1-1:0]  stream_blocks_11_attention_equery_bias;
logic                             stream_blocks_11_attention_query_bias_valid;
logic                             stream_blocks_11_attention_query_bias_ready;
logic [stream_blocks_11_attention_KEY_WEIGHT_PRECISION_0-1:0]  stream_blocks_11_attention_mkey_weight        [stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_0*stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_KEY_WEIGHT_PRECISION_1-1:0]  stream_blocks_11_attention_ekey_weight;
logic                             stream_blocks_11_attention_key_weight_valid;
logic                             stream_blocks_11_attention_key_weight_ready;
logic [stream_blocks_11_attention_KEY_BIAS_PRECISION_0-1:0]  stream_blocks_11_attention_mkey_bias        [stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_0*stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_KEY_BIAS_PRECISION_1-1:0]  stream_blocks_11_attention_ekey_bias;
logic                             stream_blocks_11_attention_key_bias_valid;
logic                             stream_blocks_11_attention_key_bias_ready;
logic [stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_0-1:0]  stream_blocks_11_attention_mvalue_weight        [stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_0*stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_1-1:0]  stream_blocks_11_attention_evalue_weight;
logic                             stream_blocks_11_attention_value_weight_valid;
logic                             stream_blocks_11_attention_value_weight_ready;
logic [stream_blocks_11_attention_VALUE_BIAS_PRECISION_0-1:0]  stream_blocks_11_attention_mvalue_bias        [stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_0*stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_VALUE_BIAS_PRECISION_1-1:0]  stream_blocks_11_attention_evalue_bias;
logic                             stream_blocks_11_attention_value_bias_valid;
logic                             stream_blocks_11_attention_value_bias_ready;
logic [stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_0-1:0]  stream_blocks_11_attention_mproj_weight        [stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_0*stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_1-1:0]  stream_blocks_11_attention_eproj_weight;
logic                             stream_blocks_11_attention_proj_weight_valid;
logic                             stream_blocks_11_attention_proj_weight_ready;
logic [stream_blocks_11_attention_PROJ_BIAS_PRECISION_0-1:0]  stream_blocks_11_attention_mproj_bias        [stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_0*stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_PROJ_BIAS_PRECISION_1-1:0]  stream_blocks_11_attention_eproj_bias;
logic                             stream_blocks_11_attention_proj_bias_valid;
logic                             stream_blocks_11_attention_proj_bias_ready;
logic [stream_blocks_11_attention_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_11_attention_mdata_out_0        [stream_blocks_11_attention_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_11_attention_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_attention_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_11_attention_edata_out_0;
logic                             stream_blocks_11_attention_data_out_0_valid;
logic                             stream_blocks_11_attention_data_out_0_ready;
// --------------------------
//   stream_blocks_11_norm2 signals
// --------------------------
logic [stream_blocks_11_norm2_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_11_norm2_mdata_in_0        [stream_blocks_11_norm2_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_11_norm2_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_norm2_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_11_norm2_edata_in_0;
logic                             stream_blocks_11_norm2_data_in_0_valid;
logic                             stream_blocks_11_norm2_data_in_0_ready;
logic [stream_blocks_11_norm2_WEIGHT_PRECISION_0-1:0]  stream_blocks_11_norm2_mweight        [stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_0*stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_norm2_WEIGHT_PRECISION_1-1:0]  stream_blocks_11_norm2_eweight;
logic                             stream_blocks_11_norm2_weight_valid;
logic                             stream_blocks_11_norm2_weight_ready;
logic [stream_blocks_11_norm2_BIAS_PRECISION_0-1:0]  stream_blocks_11_norm2_mbias        [stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_0*stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_norm2_BIAS_PRECISION_1-1:0]  stream_blocks_11_norm2_ebias;
logic                             stream_blocks_11_norm2_bias_valid;
logic                             stream_blocks_11_norm2_bias_ready;
logic [stream_blocks_11_norm2_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_11_norm2_mdata_out_0        [stream_blocks_11_norm2_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_11_norm2_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_norm2_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_11_norm2_edata_out_0;
logic                             stream_blocks_11_norm2_data_out_0_valid;
logic                             stream_blocks_11_norm2_data_out_0_ready;
// --------------------------
//   stream_blocks_11_add_1 signals
// --------------------------
logic [stream_blocks_11_add_1_DATA_IN_0_PRECISION_0-1:0]  stream_blocks_11_add_1_mdata_in_0        [stream_blocks_11_add_1_DATA_IN_0_PARALLELISM_DIM_0*stream_blocks_11_add_1_DATA_IN_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_add_1_DATA_IN_0_PRECISION_1-1:0]  stream_blocks_11_add_1_edata_in_0;
logic                             stream_blocks_11_add_1_data_in_0_valid;
logic                             stream_blocks_11_add_1_data_in_0_ready;
logic [stream_blocks_11_add_1_DATA_IN_1_PRECISION_0-1:0]  stream_blocks_11_add_1_mdata_in_1        [stream_blocks_11_add_1_DATA_IN_1_PARALLELISM_DIM_0*stream_blocks_11_add_1_DATA_IN_1_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_add_1_DATA_IN_1_PRECISION_1-1:0]  stream_blocks_11_add_1_edata_in_1;
logic                             stream_blocks_11_add_1_data_in_1_valid;
logic                             stream_blocks_11_add_1_data_in_1_ready;
logic [stream_blocks_11_add_1_DATA_OUT_0_PRECISION_0-1:0]  stream_blocks_11_add_1_mdata_out_0        [stream_blocks_11_add_1_DATA_OUT_0_PARALLELISM_DIM_0*stream_blocks_11_add_1_DATA_OUT_0_PARALLELISM_DIM_1-1:0];
logic [stream_blocks_11_add_1_DATA_OUT_0_PRECISION_1-1:0]  stream_blocks_11_add_1_edata_out_0;
logic                             stream_blocks_11_add_1_data_out_0_valid;
logic                             stream_blocks_11_add_1_data_out_0_ready;

// --------------------------
//   Component instantiation
// --------------------------

// fork2
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_mdata_in_0),
    .edata_in_0(fork2_edata_in_0),
    .data_in_0_valid(fork2_data_in_0_valid),
    .data_in_0_ready(fork2_data_in_0_ready),
        
    .mdata_out_0(fork2_mdata_out_0),
    .edata_out_0(fork2_edata_out_0),
    .data_out_0_valid(fork2_data_out_0_valid),
    .data_out_0_ready(fork2_data_out_0_ready),
        
    .mdata_out_1(fork2_mdata_out_1),
    .edata_out_1(fork2_edata_out_1),
    .data_out_1_valid(fork2_data_out_1_valid),
    .data_out_1_ready(fork2_data_out_1_ready)
);

// stream_blocks_0_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_0_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_0_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_0_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_0_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_0_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_0_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_0_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_0_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_0_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_0_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_0_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_0_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_0_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_0_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_0_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_0_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_0_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_0_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_0_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_0_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_0_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_0_linear1_mweight),
    .eweight(stream_blocks_0_linear1_eweight),
    .weight_valid(stream_blocks_0_linear1_weight_valid),
    .weight_ready(stream_blocks_0_linear1_weight_ready),
        
    .mbias(stream_blocks_0_linear1_mbias),
    .ebias(stream_blocks_0_linear1_ebias),
    .bias_valid(stream_blocks_0_linear1_bias_valid),
    .bias_ready(stream_blocks_0_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_0_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_0_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_0_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_0_linear1_data_out_0_ready)
);

stream_blocks_0_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_0_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_0_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_0_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_linear1_mweight),
    .edata_out(stream_blocks_0_linear1_eweight),
    .data_out_ready(stream_blocks_0_linear1_weight_ready),
    .data_out_valid(stream_blocks_0_linear1_weight_valid)
);

stream_blocks_0_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_0_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_0_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_0_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_0_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_linear1_mbias),
    .edata_out(stream_blocks_0_linear1_ebias),
    .data_out_ready(stream_blocks_0_linear1_bias_ready),
    .data_out_valid(stream_blocks_0_linear1_bias_valid)
);

// stream_blocks_0_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_0_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_0_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_0_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_0_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_0_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_0_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_0_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_0_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_0_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_0_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_0_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_0_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_0_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_0_act_mdata_in_0),
    .edata_in_0(stream_blocks_0_act_edata_in_0),
    .data_in_0_valid(stream_blocks_0_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_0_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_0_act_mdata_out_0),
    .edata_out_0(stream_blocks_0_act_edata_out_0),
    .data_out_0_valid(stream_blocks_0_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_0_act_data_out_0_ready)
);

// stream_blocks_0_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_0_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_0_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_0_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_0_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_0_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_0_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_0_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_0_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_0_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_0_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_0_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_0_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_0_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_0_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_0_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_0_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_0_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_0_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_0_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_0_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_0_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_0_linear2_mweight),
    .eweight(stream_blocks_0_linear2_eweight),
    .weight_valid(stream_blocks_0_linear2_weight_valid),
    .weight_ready(stream_blocks_0_linear2_weight_ready),
        
    .mbias(stream_blocks_0_linear2_mbias),
    .ebias(stream_blocks_0_linear2_ebias),
    .bias_valid(stream_blocks_0_linear2_bias_valid),
    .bias_ready(stream_blocks_0_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_0_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_0_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_0_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_0_linear2_data_out_0_ready)
);

stream_blocks_0_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_0_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_0_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_0_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_linear2_mweight),
    .edata_out(stream_blocks_0_linear2_eweight),
    .data_out_ready(stream_blocks_0_linear2_weight_ready),
    .data_out_valid(stream_blocks_0_linear2_weight_valid)
);

stream_blocks_0_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_0_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_0_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_0_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_0_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_linear2_mbias),
    .edata_out(stream_blocks_0_linear2_ebias),
    .data_out_ready(stream_blocks_0_linear2_bias_ready),
    .data_out_valid(stream_blocks_0_linear2_bias_valid)
);

// stream_blocks_0_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_0_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_0_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_0_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_0_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_0_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_0_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_0_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_0_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_0_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_0_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_0_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_0_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_0_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_0_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_0_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_0_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_0_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_0_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_0_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_0_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_0_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_0_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_0_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_0_norm1_mweight),
    .eweight(stream_blocks_0_norm1_eweight),
    .weight_valid(stream_blocks_0_norm1_weight_valid),
    .weight_ready(stream_blocks_0_norm1_weight_ready),
        
    .mbias(stream_blocks_0_norm1_mbias),
    .ebias(stream_blocks_0_norm1_ebias),
    .bias_valid(stream_blocks_0_norm1_bias_valid),
    .bias_ready(stream_blocks_0_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_0_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_0_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_0_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_0_norm1_data_out_0_ready)
);

stream_blocks_0_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_0_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_0_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_0_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_norm1_mweight),
    .edata_out(stream_blocks_0_norm1_eweight),
    .data_out_ready(stream_blocks_0_norm1_weight_ready),
    .data_out_valid(stream_blocks_0_norm1_weight_valid)
);

stream_blocks_0_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_0_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_0_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_0_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_0_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_norm1_mbias),
    .edata_out(stream_blocks_0_norm1_ebias),
    .data_out_ready(stream_blocks_0_norm1_bias_ready),
    .data_out_valid(stream_blocks_0_norm1_bias_valid)
);

// stream_blocks_0_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_0_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_0_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_0_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_0_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_0_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_0_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_0_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_0_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_0_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_0_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_0_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_0_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_0_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_0_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_0_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_0_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_0_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_0_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_0_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_0_add_mdata_in_0),
    .edata_in_0(stream_blocks_0_add_edata_in_0),
    .data_in_0_valid(stream_blocks_0_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_0_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_0_add_mdata_in_1),
    .edata_in_1(stream_blocks_0_add_edata_in_1),
    .data_in_1_valid(stream_blocks_0_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_0_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_0_add_mdata_out_0),
    .edata_out_0(stream_blocks_0_add_edata_out_0),
    .data_out_0_valid(stream_blocks_0_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_0_add_data_out_0_ready)
);

// fork2_1
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_1_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_1_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_1_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_1_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_1_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_1_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_1_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_1_mdata_in_0),
    .edata_in_0(fork2_1_edata_in_0),
    .data_in_0_valid(fork2_1_data_in_0_valid),
    .data_in_0_ready(fork2_1_data_in_0_ready),
        
    .mdata_out_0(fork2_1_mdata_out_0),
    .edata_out_0(fork2_1_edata_out_0),
    .data_out_0_valid(fork2_1_data_out_0_valid),
    .data_out_0_ready(fork2_1_data_out_0_ready),
        
    .mdata_out_1(fork2_1_mdata_out_1),
    .edata_out_1(fork2_1_edata_out_1),
    .data_out_1_valid(fork2_1_data_out_1_valid),
    .data_out_1_ready(fork2_1_data_out_1_ready)
);

// stream_blocks_0_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_0_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_0_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_0_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_0_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_0_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_0_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_0_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_0_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_0_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_0_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_0_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_0_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_0_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_0_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_0_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_0_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_0_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_0_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_0_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_0_attention_mdata_in_0),
    .edata_in_0(stream_blocks_0_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_0_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_0_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_0_attention_mquery_weight),
    .equery_weight(stream_blocks_0_attention_equery_weight),
    .query_weight_valid(stream_blocks_0_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_0_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_0_attention_mquery_bias),
    .equery_bias(stream_blocks_0_attention_equery_bias),
    .query_bias_valid(stream_blocks_0_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_0_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_0_attention_mkey_weight),
    .ekey_weight(stream_blocks_0_attention_ekey_weight),
    .key_weight_valid(stream_blocks_0_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_0_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_0_attention_mkey_bias),
    .ekey_bias(stream_blocks_0_attention_ekey_bias),
    .key_bias_valid(stream_blocks_0_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_0_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_0_attention_mvalue_weight),
    .evalue_weight(stream_blocks_0_attention_evalue_weight),
    .value_weight_valid(stream_blocks_0_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_0_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_0_attention_mvalue_bias),
    .evalue_bias(stream_blocks_0_attention_evalue_bias),
    .value_bias_valid(stream_blocks_0_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_0_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_0_attention_mproj_weight),
    .eproj_weight(stream_blocks_0_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_0_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_0_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_0_attention_mproj_bias),
    .eproj_bias(stream_blocks_0_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_0_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_0_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_0_attention_mdata_out_0),
    .edata_out_0(stream_blocks_0_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_0_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_0_attention_data_out_0_ready)
);

stream_blocks_0_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_0_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_0_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_attention_mquery_weight),
    .edata_out(stream_blocks_0_attention_equery_weight),
    .data_out_ready(stream_blocks_0_attention_query_weight_ready),
    .data_out_valid(stream_blocks_0_attention_query_weight_valid)
);

stream_blocks_0_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_0_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_0_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_0_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_0_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_attention_mquery_bias),
    .edata_out(stream_blocks_0_attention_equery_bias),
    .data_out_ready(stream_blocks_0_attention_query_bias_ready),
    .data_out_valid(stream_blocks_0_attention_query_bias_valid)
);

stream_blocks_0_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_0_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_0_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_0_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_attention_mkey_weight),
    .edata_out(stream_blocks_0_attention_ekey_weight),
    .data_out_ready(stream_blocks_0_attention_key_weight_ready),
    .data_out_valid(stream_blocks_0_attention_key_weight_valid)
);

stream_blocks_0_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_0_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_0_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_0_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_0_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_attention_mkey_bias),
    .edata_out(stream_blocks_0_attention_ekey_bias),
    .data_out_ready(stream_blocks_0_attention_key_bias_ready),
    .data_out_valid(stream_blocks_0_attention_key_bias_valid)
);

stream_blocks_0_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_0_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_0_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_attention_mvalue_weight),
    .edata_out(stream_blocks_0_attention_evalue_weight),
    .data_out_ready(stream_blocks_0_attention_value_weight_ready),
    .data_out_valid(stream_blocks_0_attention_value_weight_valid)
);

stream_blocks_0_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_0_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_0_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_0_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_0_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_attention_mvalue_bias),
    .edata_out(stream_blocks_0_attention_evalue_bias),
    .data_out_ready(stream_blocks_0_attention_value_bias_ready),
    .data_out_valid(stream_blocks_0_attention_value_bias_valid)
);

stream_blocks_0_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_0_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_0_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_attention_mproj_weight),
    .edata_out(stream_blocks_0_attention_eproj_weight),
    .data_out_ready(stream_blocks_0_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_0_attention_proj_weight_valid)
);

stream_blocks_0_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_0_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_0_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_0_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_0_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_attention_mproj_bias),
    .edata_out(stream_blocks_0_attention_eproj_bias),
    .data_out_ready(stream_blocks_0_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_0_attention_proj_bias_valid)
);

// stream_blocks_0_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_0_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_0_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_0_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_0_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_0_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_0_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_0_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_0_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_0_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_0_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_0_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_0_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_0_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_0_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_0_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_0_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_0_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_0_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_0_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_0_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_0_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_0_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_0_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_0_norm2_mweight),
    .eweight(stream_blocks_0_norm2_eweight),
    .weight_valid(stream_blocks_0_norm2_weight_valid),
    .weight_ready(stream_blocks_0_norm2_weight_ready),
        
    .mbias(stream_blocks_0_norm2_mbias),
    .ebias(stream_blocks_0_norm2_ebias),
    .bias_valid(stream_blocks_0_norm2_bias_valid),
    .bias_ready(stream_blocks_0_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_0_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_0_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_0_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_0_norm2_data_out_0_ready)
);

stream_blocks_0_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_0_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_0_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_0_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_0_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_0_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_0_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_norm2_mweight),
    .edata_out(stream_blocks_0_norm2_eweight),
    .data_out_ready(stream_blocks_0_norm2_weight_ready),
    .data_out_valid(stream_blocks_0_norm2_weight_valid)
);

stream_blocks_0_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_0_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_0_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_0_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_0_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_0_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_0_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_0_norm2_mbias),
    .edata_out(stream_blocks_0_norm2_ebias),
    .data_out_ready(stream_blocks_0_norm2_bias_ready),
    .data_out_valid(stream_blocks_0_norm2_bias_valid)
);

// stream_blocks_0_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_0_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_0_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_0_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_0_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_0_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_0_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_0_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_0_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_0_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_0_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_0_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_0_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_0_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_0_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_0_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_0_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_0_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_0_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_0_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_0_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_0_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_0_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_0_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_0_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_0_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_0_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_0_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_0_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_0_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_0_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_0_add_1_data_out_0_ready)
);

// fork2_2
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_2_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_2_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_2_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_2_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_2_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_2_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_2_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_2_mdata_in_0),
    .edata_in_0(fork2_2_edata_in_0),
    .data_in_0_valid(fork2_2_data_in_0_valid),
    .data_in_0_ready(fork2_2_data_in_0_ready),
        
    .mdata_out_0(fork2_2_mdata_out_0),
    .edata_out_0(fork2_2_edata_out_0),
    .data_out_0_valid(fork2_2_data_out_0_valid),
    .data_out_0_ready(fork2_2_data_out_0_ready),
        
    .mdata_out_1(fork2_2_mdata_out_1),
    .edata_out_1(fork2_2_edata_out_1),
    .data_out_1_valid(fork2_2_data_out_1_valid),
    .data_out_1_ready(fork2_2_data_out_1_ready)
);

// stream_blocks_1_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_1_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_1_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_1_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_1_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_1_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_1_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_1_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_1_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_1_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_1_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_1_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_1_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_1_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_1_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_1_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_1_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_1_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_1_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_1_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_1_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_1_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_1_linear1_mweight),
    .eweight(stream_blocks_1_linear1_eweight),
    .weight_valid(stream_blocks_1_linear1_weight_valid),
    .weight_ready(stream_blocks_1_linear1_weight_ready),
        
    .mbias(stream_blocks_1_linear1_mbias),
    .ebias(stream_blocks_1_linear1_ebias),
    .bias_valid(stream_blocks_1_linear1_bias_valid),
    .bias_ready(stream_blocks_1_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_1_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_1_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_1_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_1_linear1_data_out_0_ready)
);

stream_blocks_1_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_1_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_1_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_1_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_linear1_mweight),
    .edata_out(stream_blocks_1_linear1_eweight),
    .data_out_ready(stream_blocks_1_linear1_weight_ready),
    .data_out_valid(stream_blocks_1_linear1_weight_valid)
);

stream_blocks_1_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_1_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_1_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_1_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_1_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_linear1_mbias),
    .edata_out(stream_blocks_1_linear1_ebias),
    .data_out_ready(stream_blocks_1_linear1_bias_ready),
    .data_out_valid(stream_blocks_1_linear1_bias_valid)
);

// stream_blocks_1_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_1_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_1_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_1_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_1_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_1_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_1_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_1_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_1_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_1_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_1_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_1_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_1_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_1_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_1_act_mdata_in_0),
    .edata_in_0(stream_blocks_1_act_edata_in_0),
    .data_in_0_valid(stream_blocks_1_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_1_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_1_act_mdata_out_0),
    .edata_out_0(stream_blocks_1_act_edata_out_0),
    .data_out_0_valid(stream_blocks_1_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_1_act_data_out_0_ready)
);

// stream_blocks_1_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_1_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_1_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_1_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_1_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_1_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_1_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_1_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_1_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_1_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_1_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_1_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_1_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_1_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_1_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_1_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_1_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_1_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_1_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_1_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_1_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_1_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_1_linear2_mweight),
    .eweight(stream_blocks_1_linear2_eweight),
    .weight_valid(stream_blocks_1_linear2_weight_valid),
    .weight_ready(stream_blocks_1_linear2_weight_ready),
        
    .mbias(stream_blocks_1_linear2_mbias),
    .ebias(stream_blocks_1_linear2_ebias),
    .bias_valid(stream_blocks_1_linear2_bias_valid),
    .bias_ready(stream_blocks_1_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_1_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_1_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_1_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_1_linear2_data_out_0_ready)
);

stream_blocks_1_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_1_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_1_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_1_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_linear2_mweight),
    .edata_out(stream_blocks_1_linear2_eweight),
    .data_out_ready(stream_blocks_1_linear2_weight_ready),
    .data_out_valid(stream_blocks_1_linear2_weight_valid)
);

stream_blocks_1_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_1_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_1_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_1_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_1_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_linear2_mbias),
    .edata_out(stream_blocks_1_linear2_ebias),
    .data_out_ready(stream_blocks_1_linear2_bias_ready),
    .data_out_valid(stream_blocks_1_linear2_bias_valid)
);

// stream_blocks_1_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_1_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_1_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_1_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_1_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_1_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_1_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_1_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_1_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_1_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_1_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_1_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_1_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_1_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_1_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_1_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_1_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_1_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_1_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_1_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_1_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_1_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_1_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_1_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_1_norm1_mweight),
    .eweight(stream_blocks_1_norm1_eweight),
    .weight_valid(stream_blocks_1_norm1_weight_valid),
    .weight_ready(stream_blocks_1_norm1_weight_ready),
        
    .mbias(stream_blocks_1_norm1_mbias),
    .ebias(stream_blocks_1_norm1_ebias),
    .bias_valid(stream_blocks_1_norm1_bias_valid),
    .bias_ready(stream_blocks_1_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_1_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_1_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_1_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_1_norm1_data_out_0_ready)
);

stream_blocks_1_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_1_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_1_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_1_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_norm1_mweight),
    .edata_out(stream_blocks_1_norm1_eweight),
    .data_out_ready(stream_blocks_1_norm1_weight_ready),
    .data_out_valid(stream_blocks_1_norm1_weight_valid)
);

stream_blocks_1_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_1_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_1_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_1_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_1_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_norm1_mbias),
    .edata_out(stream_blocks_1_norm1_ebias),
    .data_out_ready(stream_blocks_1_norm1_bias_ready),
    .data_out_valid(stream_blocks_1_norm1_bias_valid)
);

// stream_blocks_1_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_1_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_1_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_1_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_1_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_1_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_1_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_1_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_1_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_1_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_1_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_1_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_1_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_1_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_1_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_1_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_1_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_1_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_1_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_1_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_1_add_mdata_in_0),
    .edata_in_0(stream_blocks_1_add_edata_in_0),
    .data_in_0_valid(stream_blocks_1_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_1_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_1_add_mdata_in_1),
    .edata_in_1(stream_blocks_1_add_edata_in_1),
    .data_in_1_valid(stream_blocks_1_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_1_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_1_add_mdata_out_0),
    .edata_out_0(stream_blocks_1_add_edata_out_0),
    .data_out_0_valid(stream_blocks_1_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_1_add_data_out_0_ready)
);

// fork2_3
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_3_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_3_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_3_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_3_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_3_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_3_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_3_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_3_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_3_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_3_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_3_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_3_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_3_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_3_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_3_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_3_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_3_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_3_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_3_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_3_mdata_in_0),
    .edata_in_0(fork2_3_edata_in_0),
    .data_in_0_valid(fork2_3_data_in_0_valid),
    .data_in_0_ready(fork2_3_data_in_0_ready),
        
    .mdata_out_0(fork2_3_mdata_out_0),
    .edata_out_0(fork2_3_edata_out_0),
    .data_out_0_valid(fork2_3_data_out_0_valid),
    .data_out_0_ready(fork2_3_data_out_0_ready),
        
    .mdata_out_1(fork2_3_mdata_out_1),
    .edata_out_1(fork2_3_edata_out_1),
    .data_out_1_valid(fork2_3_data_out_1_valid),
    .data_out_1_ready(fork2_3_data_out_1_ready)
);

// stream_blocks_1_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_1_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_1_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_1_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_1_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_1_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_1_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_1_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_1_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_1_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_1_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_1_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_1_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_1_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_1_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_1_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_1_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_1_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_1_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_1_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_1_attention_mdata_in_0),
    .edata_in_0(stream_blocks_1_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_1_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_1_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_1_attention_mquery_weight),
    .equery_weight(stream_blocks_1_attention_equery_weight),
    .query_weight_valid(stream_blocks_1_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_1_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_1_attention_mquery_bias),
    .equery_bias(stream_blocks_1_attention_equery_bias),
    .query_bias_valid(stream_blocks_1_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_1_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_1_attention_mkey_weight),
    .ekey_weight(stream_blocks_1_attention_ekey_weight),
    .key_weight_valid(stream_blocks_1_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_1_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_1_attention_mkey_bias),
    .ekey_bias(stream_blocks_1_attention_ekey_bias),
    .key_bias_valid(stream_blocks_1_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_1_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_1_attention_mvalue_weight),
    .evalue_weight(stream_blocks_1_attention_evalue_weight),
    .value_weight_valid(stream_blocks_1_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_1_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_1_attention_mvalue_bias),
    .evalue_bias(stream_blocks_1_attention_evalue_bias),
    .value_bias_valid(stream_blocks_1_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_1_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_1_attention_mproj_weight),
    .eproj_weight(stream_blocks_1_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_1_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_1_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_1_attention_mproj_bias),
    .eproj_bias(stream_blocks_1_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_1_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_1_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_1_attention_mdata_out_0),
    .edata_out_0(stream_blocks_1_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_1_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_1_attention_data_out_0_ready)
);

stream_blocks_1_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_1_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_1_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_attention_mquery_weight),
    .edata_out(stream_blocks_1_attention_equery_weight),
    .data_out_ready(stream_blocks_1_attention_query_weight_ready),
    .data_out_valid(stream_blocks_1_attention_query_weight_valid)
);

stream_blocks_1_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_1_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_1_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_1_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_1_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_attention_mquery_bias),
    .edata_out(stream_blocks_1_attention_equery_bias),
    .data_out_ready(stream_blocks_1_attention_query_bias_ready),
    .data_out_valid(stream_blocks_1_attention_query_bias_valid)
);

stream_blocks_1_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_1_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_1_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_1_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_attention_mkey_weight),
    .edata_out(stream_blocks_1_attention_ekey_weight),
    .data_out_ready(stream_blocks_1_attention_key_weight_ready),
    .data_out_valid(stream_blocks_1_attention_key_weight_valid)
);

stream_blocks_1_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_1_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_1_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_1_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_1_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_attention_mkey_bias),
    .edata_out(stream_blocks_1_attention_ekey_bias),
    .data_out_ready(stream_blocks_1_attention_key_bias_ready),
    .data_out_valid(stream_blocks_1_attention_key_bias_valid)
);

stream_blocks_1_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_1_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_1_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_attention_mvalue_weight),
    .edata_out(stream_blocks_1_attention_evalue_weight),
    .data_out_ready(stream_blocks_1_attention_value_weight_ready),
    .data_out_valid(stream_blocks_1_attention_value_weight_valid)
);

stream_blocks_1_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_1_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_1_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_1_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_1_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_attention_mvalue_bias),
    .edata_out(stream_blocks_1_attention_evalue_bias),
    .data_out_ready(stream_blocks_1_attention_value_bias_ready),
    .data_out_valid(stream_blocks_1_attention_value_bias_valid)
);

stream_blocks_1_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_1_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_1_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_attention_mproj_weight),
    .edata_out(stream_blocks_1_attention_eproj_weight),
    .data_out_ready(stream_blocks_1_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_1_attention_proj_weight_valid)
);

stream_blocks_1_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_1_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_1_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_1_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_1_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_attention_mproj_bias),
    .edata_out(stream_blocks_1_attention_eproj_bias),
    .data_out_ready(stream_blocks_1_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_1_attention_proj_bias_valid)
);

// stream_blocks_1_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_1_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_1_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_1_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_1_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_1_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_1_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_1_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_1_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_1_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_1_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_1_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_1_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_1_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_1_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_1_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_1_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_1_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_1_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_1_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_1_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_1_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_1_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_1_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_1_norm2_mweight),
    .eweight(stream_blocks_1_norm2_eweight),
    .weight_valid(stream_blocks_1_norm2_weight_valid),
    .weight_ready(stream_blocks_1_norm2_weight_ready),
        
    .mbias(stream_blocks_1_norm2_mbias),
    .ebias(stream_blocks_1_norm2_ebias),
    .bias_valid(stream_blocks_1_norm2_bias_valid),
    .bias_ready(stream_blocks_1_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_1_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_1_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_1_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_1_norm2_data_out_0_ready)
);

stream_blocks_1_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_1_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_1_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_1_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_1_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_1_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_1_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_norm2_mweight),
    .edata_out(stream_blocks_1_norm2_eweight),
    .data_out_ready(stream_blocks_1_norm2_weight_ready),
    .data_out_valid(stream_blocks_1_norm2_weight_valid)
);

stream_blocks_1_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_1_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_1_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_1_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_1_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_1_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_1_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_1_norm2_mbias),
    .edata_out(stream_blocks_1_norm2_ebias),
    .data_out_ready(stream_blocks_1_norm2_bias_ready),
    .data_out_valid(stream_blocks_1_norm2_bias_valid)
);

// stream_blocks_1_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_1_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_1_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_1_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_1_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_1_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_1_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_1_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_1_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_1_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_1_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_1_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_1_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_1_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_1_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_1_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_1_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_1_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_1_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_1_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_1_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_1_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_1_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_1_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_1_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_1_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_1_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_1_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_1_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_1_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_1_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_1_add_1_data_out_0_ready)
);

// fork2_4
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_4_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_4_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_4_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_4_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_4_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_4_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_4_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_4_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_4_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_4_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_4_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_4_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_4_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_4_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_4_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_4_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_4_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_4_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_4_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_4_mdata_in_0),
    .edata_in_0(fork2_4_edata_in_0),
    .data_in_0_valid(fork2_4_data_in_0_valid),
    .data_in_0_ready(fork2_4_data_in_0_ready),
        
    .mdata_out_0(fork2_4_mdata_out_0),
    .edata_out_0(fork2_4_edata_out_0),
    .data_out_0_valid(fork2_4_data_out_0_valid),
    .data_out_0_ready(fork2_4_data_out_0_ready),
        
    .mdata_out_1(fork2_4_mdata_out_1),
    .edata_out_1(fork2_4_edata_out_1),
    .data_out_1_valid(fork2_4_data_out_1_valid),
    .data_out_1_ready(fork2_4_data_out_1_ready)
);

// stream_blocks_2_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_2_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_2_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_2_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_2_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_2_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_2_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_2_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_2_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_2_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_2_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_2_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_2_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_2_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_2_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_2_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_2_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_2_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_2_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_2_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_2_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_2_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_2_linear1_mweight),
    .eweight(stream_blocks_2_linear1_eweight),
    .weight_valid(stream_blocks_2_linear1_weight_valid),
    .weight_ready(stream_blocks_2_linear1_weight_ready),
        
    .mbias(stream_blocks_2_linear1_mbias),
    .ebias(stream_blocks_2_linear1_ebias),
    .bias_valid(stream_blocks_2_linear1_bias_valid),
    .bias_ready(stream_blocks_2_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_2_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_2_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_2_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_2_linear1_data_out_0_ready)
);

stream_blocks_2_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_2_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_2_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_2_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_linear1_mweight),
    .edata_out(stream_blocks_2_linear1_eweight),
    .data_out_ready(stream_blocks_2_linear1_weight_ready),
    .data_out_valid(stream_blocks_2_linear1_weight_valid)
);

stream_blocks_2_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_2_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_2_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_2_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_2_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_linear1_mbias),
    .edata_out(stream_blocks_2_linear1_ebias),
    .data_out_ready(stream_blocks_2_linear1_bias_ready),
    .data_out_valid(stream_blocks_2_linear1_bias_valid)
);

// stream_blocks_2_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_2_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_2_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_2_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_2_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_2_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_2_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_2_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_2_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_2_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_2_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_2_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_2_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_2_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_2_act_mdata_in_0),
    .edata_in_0(stream_blocks_2_act_edata_in_0),
    .data_in_0_valid(stream_blocks_2_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_2_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_2_act_mdata_out_0),
    .edata_out_0(stream_blocks_2_act_edata_out_0),
    .data_out_0_valid(stream_blocks_2_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_2_act_data_out_0_ready)
);

// stream_blocks_2_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_2_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_2_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_2_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_2_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_2_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_2_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_2_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_2_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_2_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_2_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_2_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_2_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_2_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_2_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_2_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_2_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_2_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_2_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_2_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_2_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_2_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_2_linear2_mweight),
    .eweight(stream_blocks_2_linear2_eweight),
    .weight_valid(stream_blocks_2_linear2_weight_valid),
    .weight_ready(stream_blocks_2_linear2_weight_ready),
        
    .mbias(stream_blocks_2_linear2_mbias),
    .ebias(stream_blocks_2_linear2_ebias),
    .bias_valid(stream_blocks_2_linear2_bias_valid),
    .bias_ready(stream_blocks_2_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_2_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_2_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_2_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_2_linear2_data_out_0_ready)
);

stream_blocks_2_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_2_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_2_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_2_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_linear2_mweight),
    .edata_out(stream_blocks_2_linear2_eweight),
    .data_out_ready(stream_blocks_2_linear2_weight_ready),
    .data_out_valid(stream_blocks_2_linear2_weight_valid)
);

stream_blocks_2_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_2_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_2_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_2_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_2_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_linear2_mbias),
    .edata_out(stream_blocks_2_linear2_ebias),
    .data_out_ready(stream_blocks_2_linear2_bias_ready),
    .data_out_valid(stream_blocks_2_linear2_bias_valid)
);

// stream_blocks_2_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_2_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_2_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_2_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_2_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_2_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_2_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_2_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_2_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_2_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_2_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_2_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_2_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_2_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_2_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_2_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_2_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_2_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_2_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_2_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_2_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_2_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_2_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_2_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_2_norm1_mweight),
    .eweight(stream_blocks_2_norm1_eweight),
    .weight_valid(stream_blocks_2_norm1_weight_valid),
    .weight_ready(stream_blocks_2_norm1_weight_ready),
        
    .mbias(stream_blocks_2_norm1_mbias),
    .ebias(stream_blocks_2_norm1_ebias),
    .bias_valid(stream_blocks_2_norm1_bias_valid),
    .bias_ready(stream_blocks_2_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_2_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_2_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_2_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_2_norm1_data_out_0_ready)
);

stream_blocks_2_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_2_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_2_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_2_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_norm1_mweight),
    .edata_out(stream_blocks_2_norm1_eweight),
    .data_out_ready(stream_blocks_2_norm1_weight_ready),
    .data_out_valid(stream_blocks_2_norm1_weight_valid)
);

stream_blocks_2_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_2_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_2_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_2_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_2_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_norm1_mbias),
    .edata_out(stream_blocks_2_norm1_ebias),
    .data_out_ready(stream_blocks_2_norm1_bias_ready),
    .data_out_valid(stream_blocks_2_norm1_bias_valid)
);

// stream_blocks_2_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_2_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_2_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_2_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_2_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_2_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_2_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_2_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_2_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_2_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_2_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_2_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_2_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_2_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_2_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_2_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_2_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_2_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_2_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_2_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_2_add_mdata_in_0),
    .edata_in_0(stream_blocks_2_add_edata_in_0),
    .data_in_0_valid(stream_blocks_2_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_2_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_2_add_mdata_in_1),
    .edata_in_1(stream_blocks_2_add_edata_in_1),
    .data_in_1_valid(stream_blocks_2_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_2_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_2_add_mdata_out_0),
    .edata_out_0(stream_blocks_2_add_edata_out_0),
    .data_out_0_valid(stream_blocks_2_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_2_add_data_out_0_ready)
);

// fork2_5
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_5_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_5_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_5_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_5_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_5_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_5_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_5_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_5_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_5_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_5_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_5_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_5_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_5_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_5_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_5_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_5_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_5_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_5_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_5_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_5_mdata_in_0),
    .edata_in_0(fork2_5_edata_in_0),
    .data_in_0_valid(fork2_5_data_in_0_valid),
    .data_in_0_ready(fork2_5_data_in_0_ready),
        
    .mdata_out_0(fork2_5_mdata_out_0),
    .edata_out_0(fork2_5_edata_out_0),
    .data_out_0_valid(fork2_5_data_out_0_valid),
    .data_out_0_ready(fork2_5_data_out_0_ready),
        
    .mdata_out_1(fork2_5_mdata_out_1),
    .edata_out_1(fork2_5_edata_out_1),
    .data_out_1_valid(fork2_5_data_out_1_valid),
    .data_out_1_ready(fork2_5_data_out_1_ready)
);

// stream_blocks_2_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_2_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_2_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_2_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_2_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_2_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_2_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_2_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_2_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_2_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_2_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_2_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_2_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_2_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_2_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_2_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_2_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_2_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_2_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_2_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_2_attention_mdata_in_0),
    .edata_in_0(stream_blocks_2_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_2_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_2_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_2_attention_mquery_weight),
    .equery_weight(stream_blocks_2_attention_equery_weight),
    .query_weight_valid(stream_blocks_2_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_2_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_2_attention_mquery_bias),
    .equery_bias(stream_blocks_2_attention_equery_bias),
    .query_bias_valid(stream_blocks_2_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_2_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_2_attention_mkey_weight),
    .ekey_weight(stream_blocks_2_attention_ekey_weight),
    .key_weight_valid(stream_blocks_2_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_2_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_2_attention_mkey_bias),
    .ekey_bias(stream_blocks_2_attention_ekey_bias),
    .key_bias_valid(stream_blocks_2_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_2_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_2_attention_mvalue_weight),
    .evalue_weight(stream_blocks_2_attention_evalue_weight),
    .value_weight_valid(stream_blocks_2_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_2_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_2_attention_mvalue_bias),
    .evalue_bias(stream_blocks_2_attention_evalue_bias),
    .value_bias_valid(stream_blocks_2_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_2_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_2_attention_mproj_weight),
    .eproj_weight(stream_blocks_2_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_2_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_2_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_2_attention_mproj_bias),
    .eproj_bias(stream_blocks_2_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_2_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_2_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_2_attention_mdata_out_0),
    .edata_out_0(stream_blocks_2_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_2_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_2_attention_data_out_0_ready)
);

stream_blocks_2_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_2_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_2_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_attention_mquery_weight),
    .edata_out(stream_blocks_2_attention_equery_weight),
    .data_out_ready(stream_blocks_2_attention_query_weight_ready),
    .data_out_valid(stream_blocks_2_attention_query_weight_valid)
);

stream_blocks_2_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_2_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_2_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_2_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_2_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_attention_mquery_bias),
    .edata_out(stream_blocks_2_attention_equery_bias),
    .data_out_ready(stream_blocks_2_attention_query_bias_ready),
    .data_out_valid(stream_blocks_2_attention_query_bias_valid)
);

stream_blocks_2_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_2_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_2_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_2_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_attention_mkey_weight),
    .edata_out(stream_blocks_2_attention_ekey_weight),
    .data_out_ready(stream_blocks_2_attention_key_weight_ready),
    .data_out_valid(stream_blocks_2_attention_key_weight_valid)
);

stream_blocks_2_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_2_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_2_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_2_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_2_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_attention_mkey_bias),
    .edata_out(stream_blocks_2_attention_ekey_bias),
    .data_out_ready(stream_blocks_2_attention_key_bias_ready),
    .data_out_valid(stream_blocks_2_attention_key_bias_valid)
);

stream_blocks_2_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_2_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_2_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_attention_mvalue_weight),
    .edata_out(stream_blocks_2_attention_evalue_weight),
    .data_out_ready(stream_blocks_2_attention_value_weight_ready),
    .data_out_valid(stream_blocks_2_attention_value_weight_valid)
);

stream_blocks_2_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_2_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_2_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_2_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_2_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_attention_mvalue_bias),
    .edata_out(stream_blocks_2_attention_evalue_bias),
    .data_out_ready(stream_blocks_2_attention_value_bias_ready),
    .data_out_valid(stream_blocks_2_attention_value_bias_valid)
);

stream_blocks_2_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_2_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_2_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_attention_mproj_weight),
    .edata_out(stream_blocks_2_attention_eproj_weight),
    .data_out_ready(stream_blocks_2_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_2_attention_proj_weight_valid)
);

stream_blocks_2_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_2_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_2_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_2_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_2_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_attention_mproj_bias),
    .edata_out(stream_blocks_2_attention_eproj_bias),
    .data_out_ready(stream_blocks_2_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_2_attention_proj_bias_valid)
);

// stream_blocks_2_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_2_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_2_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_2_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_2_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_2_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_2_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_2_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_2_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_2_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_2_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_2_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_2_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_2_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_2_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_2_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_2_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_2_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_2_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_2_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_2_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_2_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_2_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_2_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_2_norm2_mweight),
    .eweight(stream_blocks_2_norm2_eweight),
    .weight_valid(stream_blocks_2_norm2_weight_valid),
    .weight_ready(stream_blocks_2_norm2_weight_ready),
        
    .mbias(stream_blocks_2_norm2_mbias),
    .ebias(stream_blocks_2_norm2_ebias),
    .bias_valid(stream_blocks_2_norm2_bias_valid),
    .bias_ready(stream_blocks_2_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_2_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_2_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_2_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_2_norm2_data_out_0_ready)
);

stream_blocks_2_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_2_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_2_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_2_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_2_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_2_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_2_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_norm2_mweight),
    .edata_out(stream_blocks_2_norm2_eweight),
    .data_out_ready(stream_blocks_2_norm2_weight_ready),
    .data_out_valid(stream_blocks_2_norm2_weight_valid)
);

stream_blocks_2_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_2_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_2_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_2_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_2_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_2_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_2_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_2_norm2_mbias),
    .edata_out(stream_blocks_2_norm2_ebias),
    .data_out_ready(stream_blocks_2_norm2_bias_ready),
    .data_out_valid(stream_blocks_2_norm2_bias_valid)
);

// stream_blocks_2_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_2_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_2_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_2_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_2_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_2_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_2_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_2_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_2_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_2_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_2_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_2_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_2_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_2_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_2_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_2_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_2_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_2_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_2_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_2_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_2_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_2_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_2_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_2_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_2_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_2_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_2_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_2_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_2_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_2_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_2_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_2_add_1_data_out_0_ready)
);

// fork2_6
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_6_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_6_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_6_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_6_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_6_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_6_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_6_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_6_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_6_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_6_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_6_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_6_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_6_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_6_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_6_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_6_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_6_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_6_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_6_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_6_mdata_in_0),
    .edata_in_0(fork2_6_edata_in_0),
    .data_in_0_valid(fork2_6_data_in_0_valid),
    .data_in_0_ready(fork2_6_data_in_0_ready),
        
    .mdata_out_0(fork2_6_mdata_out_0),
    .edata_out_0(fork2_6_edata_out_0),
    .data_out_0_valid(fork2_6_data_out_0_valid),
    .data_out_0_ready(fork2_6_data_out_0_ready),
        
    .mdata_out_1(fork2_6_mdata_out_1),
    .edata_out_1(fork2_6_edata_out_1),
    .data_out_1_valid(fork2_6_data_out_1_valid),
    .data_out_1_ready(fork2_6_data_out_1_ready)
);

// stream_blocks_3_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_3_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_3_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_3_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_3_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_3_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_3_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_3_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_3_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_3_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_3_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_3_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_3_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_3_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_3_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_3_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_3_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_3_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_3_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_3_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_3_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_3_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_3_linear1_mweight),
    .eweight(stream_blocks_3_linear1_eweight),
    .weight_valid(stream_blocks_3_linear1_weight_valid),
    .weight_ready(stream_blocks_3_linear1_weight_ready),
        
    .mbias(stream_blocks_3_linear1_mbias),
    .ebias(stream_blocks_3_linear1_ebias),
    .bias_valid(stream_blocks_3_linear1_bias_valid),
    .bias_ready(stream_blocks_3_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_3_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_3_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_3_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_3_linear1_data_out_0_ready)
);

stream_blocks_3_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_3_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_3_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_3_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_linear1_mweight),
    .edata_out(stream_blocks_3_linear1_eweight),
    .data_out_ready(stream_blocks_3_linear1_weight_ready),
    .data_out_valid(stream_blocks_3_linear1_weight_valid)
);

stream_blocks_3_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_3_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_3_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_3_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_3_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_linear1_mbias),
    .edata_out(stream_blocks_3_linear1_ebias),
    .data_out_ready(stream_blocks_3_linear1_bias_ready),
    .data_out_valid(stream_blocks_3_linear1_bias_valid)
);

// stream_blocks_3_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_3_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_3_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_3_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_3_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_3_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_3_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_3_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_3_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_3_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_3_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_3_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_3_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_3_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_3_act_mdata_in_0),
    .edata_in_0(stream_blocks_3_act_edata_in_0),
    .data_in_0_valid(stream_blocks_3_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_3_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_3_act_mdata_out_0),
    .edata_out_0(stream_blocks_3_act_edata_out_0),
    .data_out_0_valid(stream_blocks_3_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_3_act_data_out_0_ready)
);

// stream_blocks_3_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_3_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_3_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_3_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_3_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_3_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_3_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_3_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_3_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_3_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_3_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_3_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_3_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_3_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_3_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_3_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_3_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_3_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_3_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_3_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_3_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_3_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_3_linear2_mweight),
    .eweight(stream_blocks_3_linear2_eweight),
    .weight_valid(stream_blocks_3_linear2_weight_valid),
    .weight_ready(stream_blocks_3_linear2_weight_ready),
        
    .mbias(stream_blocks_3_linear2_mbias),
    .ebias(stream_blocks_3_linear2_ebias),
    .bias_valid(stream_blocks_3_linear2_bias_valid),
    .bias_ready(stream_blocks_3_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_3_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_3_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_3_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_3_linear2_data_out_0_ready)
);

stream_blocks_3_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_3_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_3_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_3_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_linear2_mweight),
    .edata_out(stream_blocks_3_linear2_eweight),
    .data_out_ready(stream_blocks_3_linear2_weight_ready),
    .data_out_valid(stream_blocks_3_linear2_weight_valid)
);

stream_blocks_3_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_3_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_3_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_3_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_3_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_linear2_mbias),
    .edata_out(stream_blocks_3_linear2_ebias),
    .data_out_ready(stream_blocks_3_linear2_bias_ready),
    .data_out_valid(stream_blocks_3_linear2_bias_valid)
);

// stream_blocks_3_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_3_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_3_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_3_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_3_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_3_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_3_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_3_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_3_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_3_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_3_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_3_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_3_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_3_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_3_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_3_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_3_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_3_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_3_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_3_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_3_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_3_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_3_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_3_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_3_norm1_mweight),
    .eweight(stream_blocks_3_norm1_eweight),
    .weight_valid(stream_blocks_3_norm1_weight_valid),
    .weight_ready(stream_blocks_3_norm1_weight_ready),
        
    .mbias(stream_blocks_3_norm1_mbias),
    .ebias(stream_blocks_3_norm1_ebias),
    .bias_valid(stream_blocks_3_norm1_bias_valid),
    .bias_ready(stream_blocks_3_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_3_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_3_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_3_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_3_norm1_data_out_0_ready)
);

stream_blocks_3_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_3_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_3_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_3_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_norm1_mweight),
    .edata_out(stream_blocks_3_norm1_eweight),
    .data_out_ready(stream_blocks_3_norm1_weight_ready),
    .data_out_valid(stream_blocks_3_norm1_weight_valid)
);

stream_blocks_3_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_3_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_3_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_3_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_3_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_norm1_mbias),
    .edata_out(stream_blocks_3_norm1_ebias),
    .data_out_ready(stream_blocks_3_norm1_bias_ready),
    .data_out_valid(stream_blocks_3_norm1_bias_valid)
);

// stream_blocks_3_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_3_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_3_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_3_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_3_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_3_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_3_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_3_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_3_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_3_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_3_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_3_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_3_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_3_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_3_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_3_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_3_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_3_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_3_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_3_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_3_add_mdata_in_0),
    .edata_in_0(stream_blocks_3_add_edata_in_0),
    .data_in_0_valid(stream_blocks_3_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_3_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_3_add_mdata_in_1),
    .edata_in_1(stream_blocks_3_add_edata_in_1),
    .data_in_1_valid(stream_blocks_3_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_3_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_3_add_mdata_out_0),
    .edata_out_0(stream_blocks_3_add_edata_out_0),
    .data_out_0_valid(stream_blocks_3_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_3_add_data_out_0_ready)
);

// fork2_7
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_7_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_7_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_7_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_7_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_7_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_7_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_7_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_7_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_7_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_7_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_7_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_7_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_7_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_7_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_7_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_7_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_7_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_7_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_7_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_7_mdata_in_0),
    .edata_in_0(fork2_7_edata_in_0),
    .data_in_0_valid(fork2_7_data_in_0_valid),
    .data_in_0_ready(fork2_7_data_in_0_ready),
        
    .mdata_out_0(fork2_7_mdata_out_0),
    .edata_out_0(fork2_7_edata_out_0),
    .data_out_0_valid(fork2_7_data_out_0_valid),
    .data_out_0_ready(fork2_7_data_out_0_ready),
        
    .mdata_out_1(fork2_7_mdata_out_1),
    .edata_out_1(fork2_7_edata_out_1),
    .data_out_1_valid(fork2_7_data_out_1_valid),
    .data_out_1_ready(fork2_7_data_out_1_ready)
);

// stream_blocks_3_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_3_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_3_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_3_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_3_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_3_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_3_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_3_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_3_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_3_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_3_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_3_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_3_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_3_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_3_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_3_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_3_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_3_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_3_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_3_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_3_attention_mdata_in_0),
    .edata_in_0(stream_blocks_3_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_3_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_3_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_3_attention_mquery_weight),
    .equery_weight(stream_blocks_3_attention_equery_weight),
    .query_weight_valid(stream_blocks_3_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_3_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_3_attention_mquery_bias),
    .equery_bias(stream_blocks_3_attention_equery_bias),
    .query_bias_valid(stream_blocks_3_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_3_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_3_attention_mkey_weight),
    .ekey_weight(stream_blocks_3_attention_ekey_weight),
    .key_weight_valid(stream_blocks_3_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_3_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_3_attention_mkey_bias),
    .ekey_bias(stream_blocks_3_attention_ekey_bias),
    .key_bias_valid(stream_blocks_3_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_3_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_3_attention_mvalue_weight),
    .evalue_weight(stream_blocks_3_attention_evalue_weight),
    .value_weight_valid(stream_blocks_3_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_3_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_3_attention_mvalue_bias),
    .evalue_bias(stream_blocks_3_attention_evalue_bias),
    .value_bias_valid(stream_blocks_3_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_3_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_3_attention_mproj_weight),
    .eproj_weight(stream_blocks_3_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_3_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_3_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_3_attention_mproj_bias),
    .eproj_bias(stream_blocks_3_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_3_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_3_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_3_attention_mdata_out_0),
    .edata_out_0(stream_blocks_3_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_3_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_3_attention_data_out_0_ready)
);

stream_blocks_3_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_3_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_3_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_attention_mquery_weight),
    .edata_out(stream_blocks_3_attention_equery_weight),
    .data_out_ready(stream_blocks_3_attention_query_weight_ready),
    .data_out_valid(stream_blocks_3_attention_query_weight_valid)
);

stream_blocks_3_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_3_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_3_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_3_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_3_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_attention_mquery_bias),
    .edata_out(stream_blocks_3_attention_equery_bias),
    .data_out_ready(stream_blocks_3_attention_query_bias_ready),
    .data_out_valid(stream_blocks_3_attention_query_bias_valid)
);

stream_blocks_3_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_3_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_3_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_3_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_attention_mkey_weight),
    .edata_out(stream_blocks_3_attention_ekey_weight),
    .data_out_ready(stream_blocks_3_attention_key_weight_ready),
    .data_out_valid(stream_blocks_3_attention_key_weight_valid)
);

stream_blocks_3_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_3_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_3_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_3_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_3_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_attention_mkey_bias),
    .edata_out(stream_blocks_3_attention_ekey_bias),
    .data_out_ready(stream_blocks_3_attention_key_bias_ready),
    .data_out_valid(stream_blocks_3_attention_key_bias_valid)
);

stream_blocks_3_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_3_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_3_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_attention_mvalue_weight),
    .edata_out(stream_blocks_3_attention_evalue_weight),
    .data_out_ready(stream_blocks_3_attention_value_weight_ready),
    .data_out_valid(stream_blocks_3_attention_value_weight_valid)
);

stream_blocks_3_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_3_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_3_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_3_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_3_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_attention_mvalue_bias),
    .edata_out(stream_blocks_3_attention_evalue_bias),
    .data_out_ready(stream_blocks_3_attention_value_bias_ready),
    .data_out_valid(stream_blocks_3_attention_value_bias_valid)
);

stream_blocks_3_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_3_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_3_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_attention_mproj_weight),
    .edata_out(stream_blocks_3_attention_eproj_weight),
    .data_out_ready(stream_blocks_3_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_3_attention_proj_weight_valid)
);

stream_blocks_3_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_3_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_3_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_3_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_3_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_attention_mproj_bias),
    .edata_out(stream_blocks_3_attention_eproj_bias),
    .data_out_ready(stream_blocks_3_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_3_attention_proj_bias_valid)
);

// stream_blocks_3_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_3_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_3_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_3_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_3_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_3_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_3_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_3_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_3_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_3_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_3_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_3_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_3_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_3_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_3_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_3_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_3_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_3_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_3_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_3_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_3_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_3_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_3_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_3_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_3_norm2_mweight),
    .eweight(stream_blocks_3_norm2_eweight),
    .weight_valid(stream_blocks_3_norm2_weight_valid),
    .weight_ready(stream_blocks_3_norm2_weight_ready),
        
    .mbias(stream_blocks_3_norm2_mbias),
    .ebias(stream_blocks_3_norm2_ebias),
    .bias_valid(stream_blocks_3_norm2_bias_valid),
    .bias_ready(stream_blocks_3_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_3_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_3_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_3_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_3_norm2_data_out_0_ready)
);

stream_blocks_3_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_3_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_3_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_3_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_3_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_3_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_3_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_norm2_mweight),
    .edata_out(stream_blocks_3_norm2_eweight),
    .data_out_ready(stream_blocks_3_norm2_weight_ready),
    .data_out_valid(stream_blocks_3_norm2_weight_valid)
);

stream_blocks_3_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_3_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_3_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_3_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_3_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_3_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_3_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_3_norm2_mbias),
    .edata_out(stream_blocks_3_norm2_ebias),
    .data_out_ready(stream_blocks_3_norm2_bias_ready),
    .data_out_valid(stream_blocks_3_norm2_bias_valid)
);

// stream_blocks_3_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_3_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_3_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_3_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_3_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_3_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_3_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_3_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_3_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_3_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_3_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_3_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_3_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_3_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_3_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_3_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_3_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_3_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_3_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_3_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_3_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_3_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_3_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_3_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_3_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_3_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_3_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_3_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_3_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_3_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_3_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_3_add_1_data_out_0_ready)
);

// fork2_8
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_8_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_8_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_8_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_8_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_8_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_8_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_8_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_8_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_8_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_8_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_8_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_8_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_8_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_8_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_8_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_8_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_8_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_8_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_8_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_8_mdata_in_0),
    .edata_in_0(fork2_8_edata_in_0),
    .data_in_0_valid(fork2_8_data_in_0_valid),
    .data_in_0_ready(fork2_8_data_in_0_ready),
        
    .mdata_out_0(fork2_8_mdata_out_0),
    .edata_out_0(fork2_8_edata_out_0),
    .data_out_0_valid(fork2_8_data_out_0_valid),
    .data_out_0_ready(fork2_8_data_out_0_ready),
        
    .mdata_out_1(fork2_8_mdata_out_1),
    .edata_out_1(fork2_8_edata_out_1),
    .data_out_1_valid(fork2_8_data_out_1_valid),
    .data_out_1_ready(fork2_8_data_out_1_ready)
);

// stream_blocks_4_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_4_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_4_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_4_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_4_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_4_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_4_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_4_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_4_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_4_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_4_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_4_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_4_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_4_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_4_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_4_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_4_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_4_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_4_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_4_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_4_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_4_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_4_linear1_mweight),
    .eweight(stream_blocks_4_linear1_eweight),
    .weight_valid(stream_blocks_4_linear1_weight_valid),
    .weight_ready(stream_blocks_4_linear1_weight_ready),
        
    .mbias(stream_blocks_4_linear1_mbias),
    .ebias(stream_blocks_4_linear1_ebias),
    .bias_valid(stream_blocks_4_linear1_bias_valid),
    .bias_ready(stream_blocks_4_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_4_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_4_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_4_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_4_linear1_data_out_0_ready)
);

stream_blocks_4_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_4_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_4_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_4_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_linear1_mweight),
    .edata_out(stream_blocks_4_linear1_eweight),
    .data_out_ready(stream_blocks_4_linear1_weight_ready),
    .data_out_valid(stream_blocks_4_linear1_weight_valid)
);

stream_blocks_4_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_4_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_4_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_4_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_4_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_linear1_mbias),
    .edata_out(stream_blocks_4_linear1_ebias),
    .data_out_ready(stream_blocks_4_linear1_bias_ready),
    .data_out_valid(stream_blocks_4_linear1_bias_valid)
);

// stream_blocks_4_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_4_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_4_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_4_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_4_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_4_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_4_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_4_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_4_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_4_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_4_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_4_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_4_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_4_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_4_act_mdata_in_0),
    .edata_in_0(stream_blocks_4_act_edata_in_0),
    .data_in_0_valid(stream_blocks_4_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_4_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_4_act_mdata_out_0),
    .edata_out_0(stream_blocks_4_act_edata_out_0),
    .data_out_0_valid(stream_blocks_4_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_4_act_data_out_0_ready)
);

// stream_blocks_4_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_4_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_4_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_4_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_4_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_4_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_4_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_4_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_4_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_4_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_4_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_4_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_4_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_4_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_4_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_4_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_4_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_4_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_4_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_4_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_4_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_4_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_4_linear2_mweight),
    .eweight(stream_blocks_4_linear2_eweight),
    .weight_valid(stream_blocks_4_linear2_weight_valid),
    .weight_ready(stream_blocks_4_linear2_weight_ready),
        
    .mbias(stream_blocks_4_linear2_mbias),
    .ebias(stream_blocks_4_linear2_ebias),
    .bias_valid(stream_blocks_4_linear2_bias_valid),
    .bias_ready(stream_blocks_4_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_4_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_4_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_4_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_4_linear2_data_out_0_ready)
);

stream_blocks_4_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_4_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_4_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_4_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_linear2_mweight),
    .edata_out(stream_blocks_4_linear2_eweight),
    .data_out_ready(stream_blocks_4_linear2_weight_ready),
    .data_out_valid(stream_blocks_4_linear2_weight_valid)
);

stream_blocks_4_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_4_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_4_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_4_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_4_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_linear2_mbias),
    .edata_out(stream_blocks_4_linear2_ebias),
    .data_out_ready(stream_blocks_4_linear2_bias_ready),
    .data_out_valid(stream_blocks_4_linear2_bias_valid)
);

// stream_blocks_4_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_4_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_4_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_4_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_4_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_4_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_4_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_4_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_4_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_4_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_4_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_4_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_4_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_4_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_4_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_4_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_4_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_4_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_4_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_4_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_4_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_4_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_4_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_4_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_4_norm1_mweight),
    .eweight(stream_blocks_4_norm1_eweight),
    .weight_valid(stream_blocks_4_norm1_weight_valid),
    .weight_ready(stream_blocks_4_norm1_weight_ready),
        
    .mbias(stream_blocks_4_norm1_mbias),
    .ebias(stream_blocks_4_norm1_ebias),
    .bias_valid(stream_blocks_4_norm1_bias_valid),
    .bias_ready(stream_blocks_4_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_4_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_4_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_4_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_4_norm1_data_out_0_ready)
);

stream_blocks_4_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_4_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_4_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_4_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_norm1_mweight),
    .edata_out(stream_blocks_4_norm1_eweight),
    .data_out_ready(stream_blocks_4_norm1_weight_ready),
    .data_out_valid(stream_blocks_4_norm1_weight_valid)
);

stream_blocks_4_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_4_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_4_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_4_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_4_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_norm1_mbias),
    .edata_out(stream_blocks_4_norm1_ebias),
    .data_out_ready(stream_blocks_4_norm1_bias_ready),
    .data_out_valid(stream_blocks_4_norm1_bias_valid)
);

// stream_blocks_4_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_4_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_4_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_4_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_4_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_4_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_4_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_4_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_4_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_4_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_4_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_4_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_4_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_4_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_4_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_4_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_4_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_4_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_4_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_4_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_4_add_mdata_in_0),
    .edata_in_0(stream_blocks_4_add_edata_in_0),
    .data_in_0_valid(stream_blocks_4_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_4_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_4_add_mdata_in_1),
    .edata_in_1(stream_blocks_4_add_edata_in_1),
    .data_in_1_valid(stream_blocks_4_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_4_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_4_add_mdata_out_0),
    .edata_out_0(stream_blocks_4_add_edata_out_0),
    .data_out_0_valid(stream_blocks_4_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_4_add_data_out_0_ready)
);

// fork2_9
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_9_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_9_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_9_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_9_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_9_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_9_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_9_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_9_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_9_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_9_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_9_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_9_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_9_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_9_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_9_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_9_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_9_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_9_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_9_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_9_mdata_in_0),
    .edata_in_0(fork2_9_edata_in_0),
    .data_in_0_valid(fork2_9_data_in_0_valid),
    .data_in_0_ready(fork2_9_data_in_0_ready),
        
    .mdata_out_0(fork2_9_mdata_out_0),
    .edata_out_0(fork2_9_edata_out_0),
    .data_out_0_valid(fork2_9_data_out_0_valid),
    .data_out_0_ready(fork2_9_data_out_0_ready),
        
    .mdata_out_1(fork2_9_mdata_out_1),
    .edata_out_1(fork2_9_edata_out_1),
    .data_out_1_valid(fork2_9_data_out_1_valid),
    .data_out_1_ready(fork2_9_data_out_1_ready)
);

// stream_blocks_4_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_4_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_4_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_4_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_4_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_4_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_4_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_4_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_4_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_4_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_4_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_4_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_4_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_4_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_4_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_4_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_4_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_4_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_4_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_4_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_4_attention_mdata_in_0),
    .edata_in_0(stream_blocks_4_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_4_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_4_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_4_attention_mquery_weight),
    .equery_weight(stream_blocks_4_attention_equery_weight),
    .query_weight_valid(stream_blocks_4_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_4_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_4_attention_mquery_bias),
    .equery_bias(stream_blocks_4_attention_equery_bias),
    .query_bias_valid(stream_blocks_4_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_4_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_4_attention_mkey_weight),
    .ekey_weight(stream_blocks_4_attention_ekey_weight),
    .key_weight_valid(stream_blocks_4_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_4_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_4_attention_mkey_bias),
    .ekey_bias(stream_blocks_4_attention_ekey_bias),
    .key_bias_valid(stream_blocks_4_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_4_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_4_attention_mvalue_weight),
    .evalue_weight(stream_blocks_4_attention_evalue_weight),
    .value_weight_valid(stream_blocks_4_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_4_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_4_attention_mvalue_bias),
    .evalue_bias(stream_blocks_4_attention_evalue_bias),
    .value_bias_valid(stream_blocks_4_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_4_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_4_attention_mproj_weight),
    .eproj_weight(stream_blocks_4_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_4_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_4_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_4_attention_mproj_bias),
    .eproj_bias(stream_blocks_4_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_4_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_4_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_4_attention_mdata_out_0),
    .edata_out_0(stream_blocks_4_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_4_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_4_attention_data_out_0_ready)
);

stream_blocks_4_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_4_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_4_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_attention_mquery_weight),
    .edata_out(stream_blocks_4_attention_equery_weight),
    .data_out_ready(stream_blocks_4_attention_query_weight_ready),
    .data_out_valid(stream_blocks_4_attention_query_weight_valid)
);

stream_blocks_4_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_4_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_4_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_4_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_4_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_attention_mquery_bias),
    .edata_out(stream_blocks_4_attention_equery_bias),
    .data_out_ready(stream_blocks_4_attention_query_bias_ready),
    .data_out_valid(stream_blocks_4_attention_query_bias_valid)
);

stream_blocks_4_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_4_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_4_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_4_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_attention_mkey_weight),
    .edata_out(stream_blocks_4_attention_ekey_weight),
    .data_out_ready(stream_blocks_4_attention_key_weight_ready),
    .data_out_valid(stream_blocks_4_attention_key_weight_valid)
);

stream_blocks_4_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_4_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_4_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_4_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_4_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_attention_mkey_bias),
    .edata_out(stream_blocks_4_attention_ekey_bias),
    .data_out_ready(stream_blocks_4_attention_key_bias_ready),
    .data_out_valid(stream_blocks_4_attention_key_bias_valid)
);

stream_blocks_4_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_4_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_4_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_attention_mvalue_weight),
    .edata_out(stream_blocks_4_attention_evalue_weight),
    .data_out_ready(stream_blocks_4_attention_value_weight_ready),
    .data_out_valid(stream_blocks_4_attention_value_weight_valid)
);

stream_blocks_4_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_4_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_4_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_4_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_4_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_attention_mvalue_bias),
    .edata_out(stream_blocks_4_attention_evalue_bias),
    .data_out_ready(stream_blocks_4_attention_value_bias_ready),
    .data_out_valid(stream_blocks_4_attention_value_bias_valid)
);

stream_blocks_4_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_4_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_4_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_attention_mproj_weight),
    .edata_out(stream_blocks_4_attention_eproj_weight),
    .data_out_ready(stream_blocks_4_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_4_attention_proj_weight_valid)
);

stream_blocks_4_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_4_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_4_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_4_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_4_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_attention_mproj_bias),
    .edata_out(stream_blocks_4_attention_eproj_bias),
    .data_out_ready(stream_blocks_4_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_4_attention_proj_bias_valid)
);

// stream_blocks_4_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_4_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_4_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_4_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_4_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_4_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_4_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_4_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_4_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_4_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_4_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_4_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_4_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_4_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_4_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_4_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_4_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_4_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_4_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_4_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_4_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_4_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_4_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_4_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_4_norm2_mweight),
    .eweight(stream_blocks_4_norm2_eweight),
    .weight_valid(stream_blocks_4_norm2_weight_valid),
    .weight_ready(stream_blocks_4_norm2_weight_ready),
        
    .mbias(stream_blocks_4_norm2_mbias),
    .ebias(stream_blocks_4_norm2_ebias),
    .bias_valid(stream_blocks_4_norm2_bias_valid),
    .bias_ready(stream_blocks_4_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_4_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_4_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_4_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_4_norm2_data_out_0_ready)
);

stream_blocks_4_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_4_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_4_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_4_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_4_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_4_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_4_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_norm2_mweight),
    .edata_out(stream_blocks_4_norm2_eweight),
    .data_out_ready(stream_blocks_4_norm2_weight_ready),
    .data_out_valid(stream_blocks_4_norm2_weight_valid)
);

stream_blocks_4_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_4_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_4_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_4_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_4_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_4_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_4_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_4_norm2_mbias),
    .edata_out(stream_blocks_4_norm2_ebias),
    .data_out_ready(stream_blocks_4_norm2_bias_ready),
    .data_out_valid(stream_blocks_4_norm2_bias_valid)
);

// stream_blocks_4_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_4_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_4_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_4_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_4_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_4_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_4_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_4_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_4_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_4_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_4_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_4_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_4_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_4_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_4_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_4_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_4_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_4_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_4_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_4_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_4_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_4_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_4_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_4_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_4_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_4_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_4_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_4_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_4_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_4_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_4_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_4_add_1_data_out_0_ready)
);

// fork2_10
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_10_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_10_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_10_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_10_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_10_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_10_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_10_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_10_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_10_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_10_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_10_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_10_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_10_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_10_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_10_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_10_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_10_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_10_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_10_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_10_mdata_in_0),
    .edata_in_0(fork2_10_edata_in_0),
    .data_in_0_valid(fork2_10_data_in_0_valid),
    .data_in_0_ready(fork2_10_data_in_0_ready),
        
    .mdata_out_0(fork2_10_mdata_out_0),
    .edata_out_0(fork2_10_edata_out_0),
    .data_out_0_valid(fork2_10_data_out_0_valid),
    .data_out_0_ready(fork2_10_data_out_0_ready),
        
    .mdata_out_1(fork2_10_mdata_out_1),
    .edata_out_1(fork2_10_edata_out_1),
    .data_out_1_valid(fork2_10_data_out_1_valid),
    .data_out_1_ready(fork2_10_data_out_1_ready)
);

// stream_blocks_5_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_5_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_5_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_5_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_5_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_5_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_5_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_5_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_5_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_5_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_5_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_5_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_5_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_5_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_5_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_5_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_5_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_5_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_5_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_5_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_5_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_5_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_5_linear1_mweight),
    .eweight(stream_blocks_5_linear1_eweight),
    .weight_valid(stream_blocks_5_linear1_weight_valid),
    .weight_ready(stream_blocks_5_linear1_weight_ready),
        
    .mbias(stream_blocks_5_linear1_mbias),
    .ebias(stream_blocks_5_linear1_ebias),
    .bias_valid(stream_blocks_5_linear1_bias_valid),
    .bias_ready(stream_blocks_5_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_5_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_5_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_5_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_5_linear1_data_out_0_ready)
);

stream_blocks_5_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_5_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_5_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_5_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_linear1_mweight),
    .edata_out(stream_blocks_5_linear1_eweight),
    .data_out_ready(stream_blocks_5_linear1_weight_ready),
    .data_out_valid(stream_blocks_5_linear1_weight_valid)
);

stream_blocks_5_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_5_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_5_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_5_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_5_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_linear1_mbias),
    .edata_out(stream_blocks_5_linear1_ebias),
    .data_out_ready(stream_blocks_5_linear1_bias_ready),
    .data_out_valid(stream_blocks_5_linear1_bias_valid)
);

// stream_blocks_5_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_5_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_5_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_5_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_5_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_5_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_5_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_5_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_5_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_5_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_5_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_5_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_5_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_5_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_5_act_mdata_in_0),
    .edata_in_0(stream_blocks_5_act_edata_in_0),
    .data_in_0_valid(stream_blocks_5_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_5_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_5_act_mdata_out_0),
    .edata_out_0(stream_blocks_5_act_edata_out_0),
    .data_out_0_valid(stream_blocks_5_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_5_act_data_out_0_ready)
);

// stream_blocks_5_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_5_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_5_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_5_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_5_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_5_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_5_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_5_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_5_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_5_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_5_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_5_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_5_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_5_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_5_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_5_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_5_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_5_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_5_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_5_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_5_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_5_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_5_linear2_mweight),
    .eweight(stream_blocks_5_linear2_eweight),
    .weight_valid(stream_blocks_5_linear2_weight_valid),
    .weight_ready(stream_blocks_5_linear2_weight_ready),
        
    .mbias(stream_blocks_5_linear2_mbias),
    .ebias(stream_blocks_5_linear2_ebias),
    .bias_valid(stream_blocks_5_linear2_bias_valid),
    .bias_ready(stream_blocks_5_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_5_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_5_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_5_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_5_linear2_data_out_0_ready)
);

stream_blocks_5_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_5_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_5_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_5_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_linear2_mweight),
    .edata_out(stream_blocks_5_linear2_eweight),
    .data_out_ready(stream_blocks_5_linear2_weight_ready),
    .data_out_valid(stream_blocks_5_linear2_weight_valid)
);

stream_blocks_5_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_5_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_5_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_5_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_5_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_linear2_mbias),
    .edata_out(stream_blocks_5_linear2_ebias),
    .data_out_ready(stream_blocks_5_linear2_bias_ready),
    .data_out_valid(stream_blocks_5_linear2_bias_valid)
);

// stream_blocks_5_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_5_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_5_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_5_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_5_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_5_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_5_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_5_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_5_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_5_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_5_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_5_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_5_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_5_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_5_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_5_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_5_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_5_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_5_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_5_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_5_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_5_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_5_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_5_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_5_norm1_mweight),
    .eweight(stream_blocks_5_norm1_eweight),
    .weight_valid(stream_blocks_5_norm1_weight_valid),
    .weight_ready(stream_blocks_5_norm1_weight_ready),
        
    .mbias(stream_blocks_5_norm1_mbias),
    .ebias(stream_blocks_5_norm1_ebias),
    .bias_valid(stream_blocks_5_norm1_bias_valid),
    .bias_ready(stream_blocks_5_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_5_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_5_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_5_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_5_norm1_data_out_0_ready)
);

stream_blocks_5_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_5_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_5_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_5_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_norm1_mweight),
    .edata_out(stream_blocks_5_norm1_eweight),
    .data_out_ready(stream_blocks_5_norm1_weight_ready),
    .data_out_valid(stream_blocks_5_norm1_weight_valid)
);

stream_blocks_5_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_5_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_5_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_5_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_5_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_norm1_mbias),
    .edata_out(stream_blocks_5_norm1_ebias),
    .data_out_ready(stream_blocks_5_norm1_bias_ready),
    .data_out_valid(stream_blocks_5_norm1_bias_valid)
);

// stream_blocks_5_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_5_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_5_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_5_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_5_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_5_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_5_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_5_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_5_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_5_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_5_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_5_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_5_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_5_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_5_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_5_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_5_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_5_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_5_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_5_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_5_add_mdata_in_0),
    .edata_in_0(stream_blocks_5_add_edata_in_0),
    .data_in_0_valid(stream_blocks_5_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_5_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_5_add_mdata_in_1),
    .edata_in_1(stream_blocks_5_add_edata_in_1),
    .data_in_1_valid(stream_blocks_5_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_5_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_5_add_mdata_out_0),
    .edata_out_0(stream_blocks_5_add_edata_out_0),
    .data_out_0_valid(stream_blocks_5_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_5_add_data_out_0_ready)
);

// fork2_11
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_11_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_11_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_11_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_11_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_11_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_11_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_11_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_11_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_11_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_11_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_11_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_11_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_11_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_11_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_11_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_11_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_11_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_11_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_11_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_11_mdata_in_0),
    .edata_in_0(fork2_11_edata_in_0),
    .data_in_0_valid(fork2_11_data_in_0_valid),
    .data_in_0_ready(fork2_11_data_in_0_ready),
        
    .mdata_out_0(fork2_11_mdata_out_0),
    .edata_out_0(fork2_11_edata_out_0),
    .data_out_0_valid(fork2_11_data_out_0_valid),
    .data_out_0_ready(fork2_11_data_out_0_ready),
        
    .mdata_out_1(fork2_11_mdata_out_1),
    .edata_out_1(fork2_11_edata_out_1),
    .data_out_1_valid(fork2_11_data_out_1_valid),
    .data_out_1_ready(fork2_11_data_out_1_ready)
);

// stream_blocks_5_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_5_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_5_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_5_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_5_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_5_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_5_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_5_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_5_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_5_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_5_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_5_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_5_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_5_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_5_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_5_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_5_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_5_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_5_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_5_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_5_attention_mdata_in_0),
    .edata_in_0(stream_blocks_5_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_5_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_5_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_5_attention_mquery_weight),
    .equery_weight(stream_blocks_5_attention_equery_weight),
    .query_weight_valid(stream_blocks_5_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_5_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_5_attention_mquery_bias),
    .equery_bias(stream_blocks_5_attention_equery_bias),
    .query_bias_valid(stream_blocks_5_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_5_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_5_attention_mkey_weight),
    .ekey_weight(stream_blocks_5_attention_ekey_weight),
    .key_weight_valid(stream_blocks_5_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_5_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_5_attention_mkey_bias),
    .ekey_bias(stream_blocks_5_attention_ekey_bias),
    .key_bias_valid(stream_blocks_5_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_5_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_5_attention_mvalue_weight),
    .evalue_weight(stream_blocks_5_attention_evalue_weight),
    .value_weight_valid(stream_blocks_5_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_5_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_5_attention_mvalue_bias),
    .evalue_bias(stream_blocks_5_attention_evalue_bias),
    .value_bias_valid(stream_blocks_5_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_5_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_5_attention_mproj_weight),
    .eproj_weight(stream_blocks_5_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_5_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_5_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_5_attention_mproj_bias),
    .eproj_bias(stream_blocks_5_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_5_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_5_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_5_attention_mdata_out_0),
    .edata_out_0(stream_blocks_5_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_5_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_5_attention_data_out_0_ready)
);

stream_blocks_5_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_5_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_5_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_attention_mquery_weight),
    .edata_out(stream_blocks_5_attention_equery_weight),
    .data_out_ready(stream_blocks_5_attention_query_weight_ready),
    .data_out_valid(stream_blocks_5_attention_query_weight_valid)
);

stream_blocks_5_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_5_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_5_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_5_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_5_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_attention_mquery_bias),
    .edata_out(stream_blocks_5_attention_equery_bias),
    .data_out_ready(stream_blocks_5_attention_query_bias_ready),
    .data_out_valid(stream_blocks_5_attention_query_bias_valid)
);

stream_blocks_5_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_5_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_5_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_5_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_attention_mkey_weight),
    .edata_out(stream_blocks_5_attention_ekey_weight),
    .data_out_ready(stream_blocks_5_attention_key_weight_ready),
    .data_out_valid(stream_blocks_5_attention_key_weight_valid)
);

stream_blocks_5_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_5_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_5_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_5_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_5_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_attention_mkey_bias),
    .edata_out(stream_blocks_5_attention_ekey_bias),
    .data_out_ready(stream_blocks_5_attention_key_bias_ready),
    .data_out_valid(stream_blocks_5_attention_key_bias_valid)
);

stream_blocks_5_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_5_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_5_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_attention_mvalue_weight),
    .edata_out(stream_blocks_5_attention_evalue_weight),
    .data_out_ready(stream_blocks_5_attention_value_weight_ready),
    .data_out_valid(stream_blocks_5_attention_value_weight_valid)
);

stream_blocks_5_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_5_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_5_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_5_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_5_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_attention_mvalue_bias),
    .edata_out(stream_blocks_5_attention_evalue_bias),
    .data_out_ready(stream_blocks_5_attention_value_bias_ready),
    .data_out_valid(stream_blocks_5_attention_value_bias_valid)
);

stream_blocks_5_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_5_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_5_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_attention_mproj_weight),
    .edata_out(stream_blocks_5_attention_eproj_weight),
    .data_out_ready(stream_blocks_5_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_5_attention_proj_weight_valid)
);

stream_blocks_5_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_5_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_5_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_5_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_5_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_attention_mproj_bias),
    .edata_out(stream_blocks_5_attention_eproj_bias),
    .data_out_ready(stream_blocks_5_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_5_attention_proj_bias_valid)
);

// stream_blocks_5_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_5_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_5_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_5_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_5_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_5_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_5_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_5_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_5_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_5_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_5_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_5_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_5_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_5_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_5_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_5_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_5_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_5_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_5_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_5_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_5_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_5_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_5_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_5_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_5_norm2_mweight),
    .eweight(stream_blocks_5_norm2_eweight),
    .weight_valid(stream_blocks_5_norm2_weight_valid),
    .weight_ready(stream_blocks_5_norm2_weight_ready),
        
    .mbias(stream_blocks_5_norm2_mbias),
    .ebias(stream_blocks_5_norm2_ebias),
    .bias_valid(stream_blocks_5_norm2_bias_valid),
    .bias_ready(stream_blocks_5_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_5_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_5_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_5_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_5_norm2_data_out_0_ready)
);

stream_blocks_5_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_5_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_5_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_5_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_5_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_5_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_5_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_norm2_mweight),
    .edata_out(stream_blocks_5_norm2_eweight),
    .data_out_ready(stream_blocks_5_norm2_weight_ready),
    .data_out_valid(stream_blocks_5_norm2_weight_valid)
);

stream_blocks_5_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_5_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_5_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_5_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_5_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_5_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_5_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_5_norm2_mbias),
    .edata_out(stream_blocks_5_norm2_ebias),
    .data_out_ready(stream_blocks_5_norm2_bias_ready),
    .data_out_valid(stream_blocks_5_norm2_bias_valid)
);

// stream_blocks_5_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_5_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_5_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_5_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_5_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_5_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_5_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_5_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_5_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_5_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_5_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_5_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_5_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_5_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_5_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_5_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_5_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_5_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_5_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_5_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_5_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_5_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_5_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_5_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_5_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_5_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_5_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_5_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_5_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_5_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_5_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_5_add_1_data_out_0_ready)
);

// fork2_12
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_12_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_12_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_12_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_12_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_12_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_12_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_12_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_12_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_12_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_12_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_12_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_12_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_12_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_12_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_12_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_12_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_12_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_12_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_12_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_12_mdata_in_0),
    .edata_in_0(fork2_12_edata_in_0),
    .data_in_0_valid(fork2_12_data_in_0_valid),
    .data_in_0_ready(fork2_12_data_in_0_ready),
        
    .mdata_out_0(fork2_12_mdata_out_0),
    .edata_out_0(fork2_12_edata_out_0),
    .data_out_0_valid(fork2_12_data_out_0_valid),
    .data_out_0_ready(fork2_12_data_out_0_ready),
        
    .mdata_out_1(fork2_12_mdata_out_1),
    .edata_out_1(fork2_12_edata_out_1),
    .data_out_1_valid(fork2_12_data_out_1_valid),
    .data_out_1_ready(fork2_12_data_out_1_ready)
);

// stream_blocks_6_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_6_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_6_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_6_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_6_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_6_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_6_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_6_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_6_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_6_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_6_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_6_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_6_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_6_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_6_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_6_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_6_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_6_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_6_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_6_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_6_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_6_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_6_linear1_mweight),
    .eweight(stream_blocks_6_linear1_eweight),
    .weight_valid(stream_blocks_6_linear1_weight_valid),
    .weight_ready(stream_blocks_6_linear1_weight_ready),
        
    .mbias(stream_blocks_6_linear1_mbias),
    .ebias(stream_blocks_6_linear1_ebias),
    .bias_valid(stream_blocks_6_linear1_bias_valid),
    .bias_ready(stream_blocks_6_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_6_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_6_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_6_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_6_linear1_data_out_0_ready)
);

stream_blocks_6_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_6_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_6_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_6_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_linear1_mweight),
    .edata_out(stream_blocks_6_linear1_eweight),
    .data_out_ready(stream_blocks_6_linear1_weight_ready),
    .data_out_valid(stream_blocks_6_linear1_weight_valid)
);

stream_blocks_6_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_6_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_6_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_6_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_6_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_linear1_mbias),
    .edata_out(stream_blocks_6_linear1_ebias),
    .data_out_ready(stream_blocks_6_linear1_bias_ready),
    .data_out_valid(stream_blocks_6_linear1_bias_valid)
);

// stream_blocks_6_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_6_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_6_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_6_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_6_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_6_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_6_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_6_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_6_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_6_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_6_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_6_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_6_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_6_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_6_act_mdata_in_0),
    .edata_in_0(stream_blocks_6_act_edata_in_0),
    .data_in_0_valid(stream_blocks_6_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_6_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_6_act_mdata_out_0),
    .edata_out_0(stream_blocks_6_act_edata_out_0),
    .data_out_0_valid(stream_blocks_6_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_6_act_data_out_0_ready)
);

// stream_blocks_6_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_6_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_6_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_6_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_6_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_6_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_6_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_6_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_6_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_6_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_6_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_6_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_6_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_6_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_6_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_6_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_6_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_6_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_6_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_6_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_6_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_6_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_6_linear2_mweight),
    .eweight(stream_blocks_6_linear2_eweight),
    .weight_valid(stream_blocks_6_linear2_weight_valid),
    .weight_ready(stream_blocks_6_linear2_weight_ready),
        
    .mbias(stream_blocks_6_linear2_mbias),
    .ebias(stream_blocks_6_linear2_ebias),
    .bias_valid(stream_blocks_6_linear2_bias_valid),
    .bias_ready(stream_blocks_6_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_6_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_6_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_6_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_6_linear2_data_out_0_ready)
);

stream_blocks_6_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_6_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_6_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_6_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_linear2_mweight),
    .edata_out(stream_blocks_6_linear2_eweight),
    .data_out_ready(stream_blocks_6_linear2_weight_ready),
    .data_out_valid(stream_blocks_6_linear2_weight_valid)
);

stream_blocks_6_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_6_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_6_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_6_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_6_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_linear2_mbias),
    .edata_out(stream_blocks_6_linear2_ebias),
    .data_out_ready(stream_blocks_6_linear2_bias_ready),
    .data_out_valid(stream_blocks_6_linear2_bias_valid)
);

// stream_blocks_6_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_6_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_6_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_6_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_6_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_6_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_6_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_6_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_6_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_6_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_6_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_6_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_6_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_6_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_6_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_6_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_6_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_6_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_6_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_6_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_6_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_6_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_6_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_6_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_6_norm1_mweight),
    .eweight(stream_blocks_6_norm1_eweight),
    .weight_valid(stream_blocks_6_norm1_weight_valid),
    .weight_ready(stream_blocks_6_norm1_weight_ready),
        
    .mbias(stream_blocks_6_norm1_mbias),
    .ebias(stream_blocks_6_norm1_ebias),
    .bias_valid(stream_blocks_6_norm1_bias_valid),
    .bias_ready(stream_blocks_6_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_6_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_6_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_6_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_6_norm1_data_out_0_ready)
);

stream_blocks_6_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_6_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_6_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_6_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_norm1_mweight),
    .edata_out(stream_blocks_6_norm1_eweight),
    .data_out_ready(stream_blocks_6_norm1_weight_ready),
    .data_out_valid(stream_blocks_6_norm1_weight_valid)
);

stream_blocks_6_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_6_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_6_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_6_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_6_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_norm1_mbias),
    .edata_out(stream_blocks_6_norm1_ebias),
    .data_out_ready(stream_blocks_6_norm1_bias_ready),
    .data_out_valid(stream_blocks_6_norm1_bias_valid)
);

// stream_blocks_6_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_6_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_6_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_6_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_6_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_6_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_6_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_6_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_6_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_6_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_6_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_6_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_6_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_6_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_6_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_6_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_6_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_6_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_6_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_6_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_6_add_mdata_in_0),
    .edata_in_0(stream_blocks_6_add_edata_in_0),
    .data_in_0_valid(stream_blocks_6_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_6_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_6_add_mdata_in_1),
    .edata_in_1(stream_blocks_6_add_edata_in_1),
    .data_in_1_valid(stream_blocks_6_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_6_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_6_add_mdata_out_0),
    .edata_out_0(stream_blocks_6_add_edata_out_0),
    .data_out_0_valid(stream_blocks_6_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_6_add_data_out_0_ready)
);

// fork2_13
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_13_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_13_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_13_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_13_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_13_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_13_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_13_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_13_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_13_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_13_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_13_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_13_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_13_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_13_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_13_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_13_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_13_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_13_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_13_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_13_mdata_in_0),
    .edata_in_0(fork2_13_edata_in_0),
    .data_in_0_valid(fork2_13_data_in_0_valid),
    .data_in_0_ready(fork2_13_data_in_0_ready),
        
    .mdata_out_0(fork2_13_mdata_out_0),
    .edata_out_0(fork2_13_edata_out_0),
    .data_out_0_valid(fork2_13_data_out_0_valid),
    .data_out_0_ready(fork2_13_data_out_0_ready),
        
    .mdata_out_1(fork2_13_mdata_out_1),
    .edata_out_1(fork2_13_edata_out_1),
    .data_out_1_valid(fork2_13_data_out_1_valid),
    .data_out_1_ready(fork2_13_data_out_1_ready)
);

// stream_blocks_6_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_6_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_6_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_6_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_6_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_6_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_6_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_6_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_6_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_6_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_6_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_6_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_6_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_6_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_6_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_6_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_6_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_6_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_6_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_6_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_6_attention_mdata_in_0),
    .edata_in_0(stream_blocks_6_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_6_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_6_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_6_attention_mquery_weight),
    .equery_weight(stream_blocks_6_attention_equery_weight),
    .query_weight_valid(stream_blocks_6_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_6_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_6_attention_mquery_bias),
    .equery_bias(stream_blocks_6_attention_equery_bias),
    .query_bias_valid(stream_blocks_6_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_6_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_6_attention_mkey_weight),
    .ekey_weight(stream_blocks_6_attention_ekey_weight),
    .key_weight_valid(stream_blocks_6_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_6_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_6_attention_mkey_bias),
    .ekey_bias(stream_blocks_6_attention_ekey_bias),
    .key_bias_valid(stream_blocks_6_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_6_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_6_attention_mvalue_weight),
    .evalue_weight(stream_blocks_6_attention_evalue_weight),
    .value_weight_valid(stream_blocks_6_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_6_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_6_attention_mvalue_bias),
    .evalue_bias(stream_blocks_6_attention_evalue_bias),
    .value_bias_valid(stream_blocks_6_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_6_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_6_attention_mproj_weight),
    .eproj_weight(stream_blocks_6_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_6_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_6_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_6_attention_mproj_bias),
    .eproj_bias(stream_blocks_6_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_6_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_6_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_6_attention_mdata_out_0),
    .edata_out_0(stream_blocks_6_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_6_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_6_attention_data_out_0_ready)
);

stream_blocks_6_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_6_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_6_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_attention_mquery_weight),
    .edata_out(stream_blocks_6_attention_equery_weight),
    .data_out_ready(stream_blocks_6_attention_query_weight_ready),
    .data_out_valid(stream_blocks_6_attention_query_weight_valid)
);

stream_blocks_6_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_6_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_6_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_6_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_6_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_attention_mquery_bias),
    .edata_out(stream_blocks_6_attention_equery_bias),
    .data_out_ready(stream_blocks_6_attention_query_bias_ready),
    .data_out_valid(stream_blocks_6_attention_query_bias_valid)
);

stream_blocks_6_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_6_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_6_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_6_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_attention_mkey_weight),
    .edata_out(stream_blocks_6_attention_ekey_weight),
    .data_out_ready(stream_blocks_6_attention_key_weight_ready),
    .data_out_valid(stream_blocks_6_attention_key_weight_valid)
);

stream_blocks_6_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_6_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_6_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_6_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_6_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_attention_mkey_bias),
    .edata_out(stream_blocks_6_attention_ekey_bias),
    .data_out_ready(stream_blocks_6_attention_key_bias_ready),
    .data_out_valid(stream_blocks_6_attention_key_bias_valid)
);

stream_blocks_6_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_6_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_6_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_attention_mvalue_weight),
    .edata_out(stream_blocks_6_attention_evalue_weight),
    .data_out_ready(stream_blocks_6_attention_value_weight_ready),
    .data_out_valid(stream_blocks_6_attention_value_weight_valid)
);

stream_blocks_6_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_6_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_6_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_6_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_6_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_attention_mvalue_bias),
    .edata_out(stream_blocks_6_attention_evalue_bias),
    .data_out_ready(stream_blocks_6_attention_value_bias_ready),
    .data_out_valid(stream_blocks_6_attention_value_bias_valid)
);

stream_blocks_6_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_6_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_6_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_attention_mproj_weight),
    .edata_out(stream_blocks_6_attention_eproj_weight),
    .data_out_ready(stream_blocks_6_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_6_attention_proj_weight_valid)
);

stream_blocks_6_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_6_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_6_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_6_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_6_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_attention_mproj_bias),
    .edata_out(stream_blocks_6_attention_eproj_bias),
    .data_out_ready(stream_blocks_6_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_6_attention_proj_bias_valid)
);

// stream_blocks_6_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_6_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_6_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_6_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_6_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_6_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_6_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_6_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_6_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_6_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_6_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_6_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_6_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_6_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_6_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_6_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_6_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_6_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_6_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_6_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_6_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_6_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_6_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_6_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_6_norm2_mweight),
    .eweight(stream_blocks_6_norm2_eweight),
    .weight_valid(stream_blocks_6_norm2_weight_valid),
    .weight_ready(stream_blocks_6_norm2_weight_ready),
        
    .mbias(stream_blocks_6_norm2_mbias),
    .ebias(stream_blocks_6_norm2_ebias),
    .bias_valid(stream_blocks_6_norm2_bias_valid),
    .bias_ready(stream_blocks_6_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_6_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_6_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_6_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_6_norm2_data_out_0_ready)
);

stream_blocks_6_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_6_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_6_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_6_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_6_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_6_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_6_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_norm2_mweight),
    .edata_out(stream_blocks_6_norm2_eweight),
    .data_out_ready(stream_blocks_6_norm2_weight_ready),
    .data_out_valid(stream_blocks_6_norm2_weight_valid)
);

stream_blocks_6_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_6_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_6_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_6_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_6_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_6_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_6_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_6_norm2_mbias),
    .edata_out(stream_blocks_6_norm2_ebias),
    .data_out_ready(stream_blocks_6_norm2_bias_ready),
    .data_out_valid(stream_blocks_6_norm2_bias_valid)
);

// stream_blocks_6_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_6_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_6_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_6_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_6_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_6_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_6_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_6_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_6_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_6_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_6_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_6_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_6_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_6_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_6_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_6_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_6_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_6_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_6_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_6_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_6_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_6_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_6_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_6_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_6_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_6_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_6_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_6_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_6_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_6_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_6_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_6_add_1_data_out_0_ready)
);

// fork2_14
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_14_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_14_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_14_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_14_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_14_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_14_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_14_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_14_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_14_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_14_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_14_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_14_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_14_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_14_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_14_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_14_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_14_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_14_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_14_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_14_mdata_in_0),
    .edata_in_0(fork2_14_edata_in_0),
    .data_in_0_valid(fork2_14_data_in_0_valid),
    .data_in_0_ready(fork2_14_data_in_0_ready),
        
    .mdata_out_0(fork2_14_mdata_out_0),
    .edata_out_0(fork2_14_edata_out_0),
    .data_out_0_valid(fork2_14_data_out_0_valid),
    .data_out_0_ready(fork2_14_data_out_0_ready),
        
    .mdata_out_1(fork2_14_mdata_out_1),
    .edata_out_1(fork2_14_edata_out_1),
    .data_out_1_valid(fork2_14_data_out_1_valid),
    .data_out_1_ready(fork2_14_data_out_1_ready)
);

// stream_blocks_7_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_7_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_7_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_7_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_7_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_7_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_7_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_7_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_7_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_7_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_7_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_7_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_7_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_7_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_7_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_7_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_7_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_7_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_7_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_7_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_7_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_7_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_7_linear1_mweight),
    .eweight(stream_blocks_7_linear1_eweight),
    .weight_valid(stream_blocks_7_linear1_weight_valid),
    .weight_ready(stream_blocks_7_linear1_weight_ready),
        
    .mbias(stream_blocks_7_linear1_mbias),
    .ebias(stream_blocks_7_linear1_ebias),
    .bias_valid(stream_blocks_7_linear1_bias_valid),
    .bias_ready(stream_blocks_7_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_7_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_7_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_7_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_7_linear1_data_out_0_ready)
);

stream_blocks_7_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_7_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_7_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_7_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_linear1_mweight),
    .edata_out(stream_blocks_7_linear1_eweight),
    .data_out_ready(stream_blocks_7_linear1_weight_ready),
    .data_out_valid(stream_blocks_7_linear1_weight_valid)
);

stream_blocks_7_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_7_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_7_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_7_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_7_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_linear1_mbias),
    .edata_out(stream_blocks_7_linear1_ebias),
    .data_out_ready(stream_blocks_7_linear1_bias_ready),
    .data_out_valid(stream_blocks_7_linear1_bias_valid)
);

// stream_blocks_7_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_7_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_7_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_7_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_7_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_7_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_7_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_7_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_7_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_7_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_7_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_7_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_7_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_7_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_7_act_mdata_in_0),
    .edata_in_0(stream_blocks_7_act_edata_in_0),
    .data_in_0_valid(stream_blocks_7_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_7_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_7_act_mdata_out_0),
    .edata_out_0(stream_blocks_7_act_edata_out_0),
    .data_out_0_valid(stream_blocks_7_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_7_act_data_out_0_ready)
);

// stream_blocks_7_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_7_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_7_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_7_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_7_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_7_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_7_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_7_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_7_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_7_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_7_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_7_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_7_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_7_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_7_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_7_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_7_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_7_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_7_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_7_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_7_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_7_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_7_linear2_mweight),
    .eweight(stream_blocks_7_linear2_eweight),
    .weight_valid(stream_blocks_7_linear2_weight_valid),
    .weight_ready(stream_blocks_7_linear2_weight_ready),
        
    .mbias(stream_blocks_7_linear2_mbias),
    .ebias(stream_blocks_7_linear2_ebias),
    .bias_valid(stream_blocks_7_linear2_bias_valid),
    .bias_ready(stream_blocks_7_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_7_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_7_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_7_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_7_linear2_data_out_0_ready)
);

stream_blocks_7_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_7_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_7_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_7_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_linear2_mweight),
    .edata_out(stream_blocks_7_linear2_eweight),
    .data_out_ready(stream_blocks_7_linear2_weight_ready),
    .data_out_valid(stream_blocks_7_linear2_weight_valid)
);

stream_blocks_7_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_7_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_7_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_7_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_7_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_linear2_mbias),
    .edata_out(stream_blocks_7_linear2_ebias),
    .data_out_ready(stream_blocks_7_linear2_bias_ready),
    .data_out_valid(stream_blocks_7_linear2_bias_valid)
);

// stream_blocks_7_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_7_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_7_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_7_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_7_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_7_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_7_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_7_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_7_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_7_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_7_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_7_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_7_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_7_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_7_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_7_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_7_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_7_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_7_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_7_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_7_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_7_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_7_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_7_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_7_norm1_mweight),
    .eweight(stream_blocks_7_norm1_eweight),
    .weight_valid(stream_blocks_7_norm1_weight_valid),
    .weight_ready(stream_blocks_7_norm1_weight_ready),
        
    .mbias(stream_blocks_7_norm1_mbias),
    .ebias(stream_blocks_7_norm1_ebias),
    .bias_valid(stream_blocks_7_norm1_bias_valid),
    .bias_ready(stream_blocks_7_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_7_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_7_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_7_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_7_norm1_data_out_0_ready)
);

stream_blocks_7_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_7_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_7_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_7_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_norm1_mweight),
    .edata_out(stream_blocks_7_norm1_eweight),
    .data_out_ready(stream_blocks_7_norm1_weight_ready),
    .data_out_valid(stream_blocks_7_norm1_weight_valid)
);

stream_blocks_7_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_7_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_7_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_7_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_7_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_norm1_mbias),
    .edata_out(stream_blocks_7_norm1_ebias),
    .data_out_ready(stream_blocks_7_norm1_bias_ready),
    .data_out_valid(stream_blocks_7_norm1_bias_valid)
);

// stream_blocks_7_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_7_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_7_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_7_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_7_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_7_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_7_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_7_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_7_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_7_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_7_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_7_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_7_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_7_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_7_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_7_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_7_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_7_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_7_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_7_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_7_add_mdata_in_0),
    .edata_in_0(stream_blocks_7_add_edata_in_0),
    .data_in_0_valid(stream_blocks_7_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_7_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_7_add_mdata_in_1),
    .edata_in_1(stream_blocks_7_add_edata_in_1),
    .data_in_1_valid(stream_blocks_7_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_7_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_7_add_mdata_out_0),
    .edata_out_0(stream_blocks_7_add_edata_out_0),
    .data_out_0_valid(stream_blocks_7_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_7_add_data_out_0_ready)
);

// fork2_15
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_15_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_15_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_15_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_15_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_15_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_15_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_15_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_15_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_15_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_15_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_15_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_15_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_15_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_15_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_15_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_15_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_15_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_15_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_15_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_15_mdata_in_0),
    .edata_in_0(fork2_15_edata_in_0),
    .data_in_0_valid(fork2_15_data_in_0_valid),
    .data_in_0_ready(fork2_15_data_in_0_ready),
        
    .mdata_out_0(fork2_15_mdata_out_0),
    .edata_out_0(fork2_15_edata_out_0),
    .data_out_0_valid(fork2_15_data_out_0_valid),
    .data_out_0_ready(fork2_15_data_out_0_ready),
        
    .mdata_out_1(fork2_15_mdata_out_1),
    .edata_out_1(fork2_15_edata_out_1),
    .data_out_1_valid(fork2_15_data_out_1_valid),
    .data_out_1_ready(fork2_15_data_out_1_ready)
);

// stream_blocks_7_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_7_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_7_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_7_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_7_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_7_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_7_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_7_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_7_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_7_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_7_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_7_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_7_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_7_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_7_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_7_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_7_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_7_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_7_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_7_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_7_attention_mdata_in_0),
    .edata_in_0(stream_blocks_7_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_7_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_7_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_7_attention_mquery_weight),
    .equery_weight(stream_blocks_7_attention_equery_weight),
    .query_weight_valid(stream_blocks_7_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_7_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_7_attention_mquery_bias),
    .equery_bias(stream_blocks_7_attention_equery_bias),
    .query_bias_valid(stream_blocks_7_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_7_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_7_attention_mkey_weight),
    .ekey_weight(stream_blocks_7_attention_ekey_weight),
    .key_weight_valid(stream_blocks_7_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_7_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_7_attention_mkey_bias),
    .ekey_bias(stream_blocks_7_attention_ekey_bias),
    .key_bias_valid(stream_blocks_7_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_7_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_7_attention_mvalue_weight),
    .evalue_weight(stream_blocks_7_attention_evalue_weight),
    .value_weight_valid(stream_blocks_7_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_7_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_7_attention_mvalue_bias),
    .evalue_bias(stream_blocks_7_attention_evalue_bias),
    .value_bias_valid(stream_blocks_7_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_7_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_7_attention_mproj_weight),
    .eproj_weight(stream_blocks_7_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_7_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_7_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_7_attention_mproj_bias),
    .eproj_bias(stream_blocks_7_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_7_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_7_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_7_attention_mdata_out_0),
    .edata_out_0(stream_blocks_7_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_7_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_7_attention_data_out_0_ready)
);

stream_blocks_7_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_7_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_7_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_attention_mquery_weight),
    .edata_out(stream_blocks_7_attention_equery_weight),
    .data_out_ready(stream_blocks_7_attention_query_weight_ready),
    .data_out_valid(stream_blocks_7_attention_query_weight_valid)
);

stream_blocks_7_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_7_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_7_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_7_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_7_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_attention_mquery_bias),
    .edata_out(stream_blocks_7_attention_equery_bias),
    .data_out_ready(stream_blocks_7_attention_query_bias_ready),
    .data_out_valid(stream_blocks_7_attention_query_bias_valid)
);

stream_blocks_7_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_7_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_7_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_7_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_attention_mkey_weight),
    .edata_out(stream_blocks_7_attention_ekey_weight),
    .data_out_ready(stream_blocks_7_attention_key_weight_ready),
    .data_out_valid(stream_blocks_7_attention_key_weight_valid)
);

stream_blocks_7_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_7_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_7_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_7_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_7_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_attention_mkey_bias),
    .edata_out(stream_blocks_7_attention_ekey_bias),
    .data_out_ready(stream_blocks_7_attention_key_bias_ready),
    .data_out_valid(stream_blocks_7_attention_key_bias_valid)
);

stream_blocks_7_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_7_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_7_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_attention_mvalue_weight),
    .edata_out(stream_blocks_7_attention_evalue_weight),
    .data_out_ready(stream_blocks_7_attention_value_weight_ready),
    .data_out_valid(stream_blocks_7_attention_value_weight_valid)
);

stream_blocks_7_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_7_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_7_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_7_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_7_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_attention_mvalue_bias),
    .edata_out(stream_blocks_7_attention_evalue_bias),
    .data_out_ready(stream_blocks_7_attention_value_bias_ready),
    .data_out_valid(stream_blocks_7_attention_value_bias_valid)
);

stream_blocks_7_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_7_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_7_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_attention_mproj_weight),
    .edata_out(stream_blocks_7_attention_eproj_weight),
    .data_out_ready(stream_blocks_7_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_7_attention_proj_weight_valid)
);

stream_blocks_7_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_7_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_7_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_7_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_7_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_attention_mproj_bias),
    .edata_out(stream_blocks_7_attention_eproj_bias),
    .data_out_ready(stream_blocks_7_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_7_attention_proj_bias_valid)
);

// stream_blocks_7_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_7_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_7_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_7_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_7_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_7_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_7_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_7_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_7_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_7_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_7_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_7_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_7_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_7_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_7_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_7_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_7_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_7_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_7_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_7_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_7_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_7_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_7_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_7_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_7_norm2_mweight),
    .eweight(stream_blocks_7_norm2_eweight),
    .weight_valid(stream_blocks_7_norm2_weight_valid),
    .weight_ready(stream_blocks_7_norm2_weight_ready),
        
    .mbias(stream_blocks_7_norm2_mbias),
    .ebias(stream_blocks_7_norm2_ebias),
    .bias_valid(stream_blocks_7_norm2_bias_valid),
    .bias_ready(stream_blocks_7_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_7_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_7_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_7_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_7_norm2_data_out_0_ready)
);

stream_blocks_7_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_7_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_7_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_7_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_7_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_7_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_7_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_norm2_mweight),
    .edata_out(stream_blocks_7_norm2_eweight),
    .data_out_ready(stream_blocks_7_norm2_weight_ready),
    .data_out_valid(stream_blocks_7_norm2_weight_valid)
);

stream_blocks_7_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_7_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_7_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_7_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_7_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_7_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_7_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_7_norm2_mbias),
    .edata_out(stream_blocks_7_norm2_ebias),
    .data_out_ready(stream_blocks_7_norm2_bias_ready),
    .data_out_valid(stream_blocks_7_norm2_bias_valid)
);

// stream_blocks_7_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_7_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_7_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_7_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_7_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_7_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_7_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_7_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_7_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_7_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_7_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_7_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_7_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_7_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_7_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_7_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_7_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_7_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_7_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_7_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_7_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_7_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_7_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_7_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_7_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_7_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_7_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_7_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_7_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_7_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_7_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_7_add_1_data_out_0_ready)
);

// fork2_16
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_16_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_16_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_16_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_16_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_16_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_16_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_16_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_16_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_16_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_16_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_16_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_16_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_16_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_16_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_16_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_16_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_16_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_16_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_16_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_16_mdata_in_0),
    .edata_in_0(fork2_16_edata_in_0),
    .data_in_0_valid(fork2_16_data_in_0_valid),
    .data_in_0_ready(fork2_16_data_in_0_ready),
        
    .mdata_out_0(fork2_16_mdata_out_0),
    .edata_out_0(fork2_16_edata_out_0),
    .data_out_0_valid(fork2_16_data_out_0_valid),
    .data_out_0_ready(fork2_16_data_out_0_ready),
        
    .mdata_out_1(fork2_16_mdata_out_1),
    .edata_out_1(fork2_16_edata_out_1),
    .data_out_1_valid(fork2_16_data_out_1_valid),
    .data_out_1_ready(fork2_16_data_out_1_ready)
);

// stream_blocks_8_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_8_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_8_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_8_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_8_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_8_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_8_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_8_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_8_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_8_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_8_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_8_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_8_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_8_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_8_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_8_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_8_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_8_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_8_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_8_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_8_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_8_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_8_linear1_mweight),
    .eweight(stream_blocks_8_linear1_eweight),
    .weight_valid(stream_blocks_8_linear1_weight_valid),
    .weight_ready(stream_blocks_8_linear1_weight_ready),
        
    .mbias(stream_blocks_8_linear1_mbias),
    .ebias(stream_blocks_8_linear1_ebias),
    .bias_valid(stream_blocks_8_linear1_bias_valid),
    .bias_ready(stream_blocks_8_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_8_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_8_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_8_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_8_linear1_data_out_0_ready)
);

stream_blocks_8_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_8_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_8_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_8_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_linear1_mweight),
    .edata_out(stream_blocks_8_linear1_eweight),
    .data_out_ready(stream_blocks_8_linear1_weight_ready),
    .data_out_valid(stream_blocks_8_linear1_weight_valid)
);

stream_blocks_8_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_8_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_8_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_8_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_8_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_linear1_mbias),
    .edata_out(stream_blocks_8_linear1_ebias),
    .data_out_ready(stream_blocks_8_linear1_bias_ready),
    .data_out_valid(stream_blocks_8_linear1_bias_valid)
);

// stream_blocks_8_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_8_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_8_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_8_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_8_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_8_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_8_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_8_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_8_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_8_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_8_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_8_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_8_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_8_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_8_act_mdata_in_0),
    .edata_in_0(stream_blocks_8_act_edata_in_0),
    .data_in_0_valid(stream_blocks_8_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_8_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_8_act_mdata_out_0),
    .edata_out_0(stream_blocks_8_act_edata_out_0),
    .data_out_0_valid(stream_blocks_8_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_8_act_data_out_0_ready)
);

// stream_blocks_8_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_8_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_8_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_8_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_8_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_8_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_8_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_8_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_8_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_8_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_8_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_8_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_8_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_8_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_8_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_8_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_8_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_8_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_8_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_8_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_8_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_8_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_8_linear2_mweight),
    .eweight(stream_blocks_8_linear2_eweight),
    .weight_valid(stream_blocks_8_linear2_weight_valid),
    .weight_ready(stream_blocks_8_linear2_weight_ready),
        
    .mbias(stream_blocks_8_linear2_mbias),
    .ebias(stream_blocks_8_linear2_ebias),
    .bias_valid(stream_blocks_8_linear2_bias_valid),
    .bias_ready(stream_blocks_8_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_8_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_8_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_8_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_8_linear2_data_out_0_ready)
);

stream_blocks_8_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_8_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_8_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_8_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_linear2_mweight),
    .edata_out(stream_blocks_8_linear2_eweight),
    .data_out_ready(stream_blocks_8_linear2_weight_ready),
    .data_out_valid(stream_blocks_8_linear2_weight_valid)
);

stream_blocks_8_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_8_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_8_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_8_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_8_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_linear2_mbias),
    .edata_out(stream_blocks_8_linear2_ebias),
    .data_out_ready(stream_blocks_8_linear2_bias_ready),
    .data_out_valid(stream_blocks_8_linear2_bias_valid)
);

// stream_blocks_8_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_8_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_8_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_8_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_8_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_8_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_8_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_8_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_8_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_8_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_8_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_8_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_8_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_8_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_8_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_8_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_8_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_8_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_8_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_8_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_8_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_8_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_8_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_8_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_8_norm1_mweight),
    .eweight(stream_blocks_8_norm1_eweight),
    .weight_valid(stream_blocks_8_norm1_weight_valid),
    .weight_ready(stream_blocks_8_norm1_weight_ready),
        
    .mbias(stream_blocks_8_norm1_mbias),
    .ebias(stream_blocks_8_norm1_ebias),
    .bias_valid(stream_blocks_8_norm1_bias_valid),
    .bias_ready(stream_blocks_8_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_8_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_8_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_8_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_8_norm1_data_out_0_ready)
);

stream_blocks_8_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_8_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_8_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_8_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_norm1_mweight),
    .edata_out(stream_blocks_8_norm1_eweight),
    .data_out_ready(stream_blocks_8_norm1_weight_ready),
    .data_out_valid(stream_blocks_8_norm1_weight_valid)
);

stream_blocks_8_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_8_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_8_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_8_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_8_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_norm1_mbias),
    .edata_out(stream_blocks_8_norm1_ebias),
    .data_out_ready(stream_blocks_8_norm1_bias_ready),
    .data_out_valid(stream_blocks_8_norm1_bias_valid)
);

// stream_blocks_8_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_8_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_8_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_8_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_8_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_8_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_8_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_8_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_8_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_8_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_8_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_8_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_8_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_8_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_8_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_8_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_8_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_8_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_8_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_8_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_8_add_mdata_in_0),
    .edata_in_0(stream_blocks_8_add_edata_in_0),
    .data_in_0_valid(stream_blocks_8_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_8_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_8_add_mdata_in_1),
    .edata_in_1(stream_blocks_8_add_edata_in_1),
    .data_in_1_valid(stream_blocks_8_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_8_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_8_add_mdata_out_0),
    .edata_out_0(stream_blocks_8_add_edata_out_0),
    .data_out_0_valid(stream_blocks_8_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_8_add_data_out_0_ready)
);

// fork2_17
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_17_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_17_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_17_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_17_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_17_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_17_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_17_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_17_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_17_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_17_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_17_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_17_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_17_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_17_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_17_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_17_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_17_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_17_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_17_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_17_mdata_in_0),
    .edata_in_0(fork2_17_edata_in_0),
    .data_in_0_valid(fork2_17_data_in_0_valid),
    .data_in_0_ready(fork2_17_data_in_0_ready),
        
    .mdata_out_0(fork2_17_mdata_out_0),
    .edata_out_0(fork2_17_edata_out_0),
    .data_out_0_valid(fork2_17_data_out_0_valid),
    .data_out_0_ready(fork2_17_data_out_0_ready),
        
    .mdata_out_1(fork2_17_mdata_out_1),
    .edata_out_1(fork2_17_edata_out_1),
    .data_out_1_valid(fork2_17_data_out_1_valid),
    .data_out_1_ready(fork2_17_data_out_1_ready)
);

// stream_blocks_8_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_8_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_8_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_8_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_8_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_8_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_8_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_8_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_8_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_8_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_8_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_8_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_8_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_8_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_8_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_8_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_8_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_8_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_8_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_8_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_8_attention_mdata_in_0),
    .edata_in_0(stream_blocks_8_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_8_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_8_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_8_attention_mquery_weight),
    .equery_weight(stream_blocks_8_attention_equery_weight),
    .query_weight_valid(stream_blocks_8_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_8_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_8_attention_mquery_bias),
    .equery_bias(stream_blocks_8_attention_equery_bias),
    .query_bias_valid(stream_blocks_8_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_8_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_8_attention_mkey_weight),
    .ekey_weight(stream_blocks_8_attention_ekey_weight),
    .key_weight_valid(stream_blocks_8_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_8_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_8_attention_mkey_bias),
    .ekey_bias(stream_blocks_8_attention_ekey_bias),
    .key_bias_valid(stream_blocks_8_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_8_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_8_attention_mvalue_weight),
    .evalue_weight(stream_blocks_8_attention_evalue_weight),
    .value_weight_valid(stream_blocks_8_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_8_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_8_attention_mvalue_bias),
    .evalue_bias(stream_blocks_8_attention_evalue_bias),
    .value_bias_valid(stream_blocks_8_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_8_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_8_attention_mproj_weight),
    .eproj_weight(stream_blocks_8_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_8_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_8_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_8_attention_mproj_bias),
    .eproj_bias(stream_blocks_8_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_8_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_8_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_8_attention_mdata_out_0),
    .edata_out_0(stream_blocks_8_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_8_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_8_attention_data_out_0_ready)
);

stream_blocks_8_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_8_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_8_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_attention_mquery_weight),
    .edata_out(stream_blocks_8_attention_equery_weight),
    .data_out_ready(stream_blocks_8_attention_query_weight_ready),
    .data_out_valid(stream_blocks_8_attention_query_weight_valid)
);

stream_blocks_8_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_8_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_8_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_8_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_8_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_attention_mquery_bias),
    .edata_out(stream_blocks_8_attention_equery_bias),
    .data_out_ready(stream_blocks_8_attention_query_bias_ready),
    .data_out_valid(stream_blocks_8_attention_query_bias_valid)
);

stream_blocks_8_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_8_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_8_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_8_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_attention_mkey_weight),
    .edata_out(stream_blocks_8_attention_ekey_weight),
    .data_out_ready(stream_blocks_8_attention_key_weight_ready),
    .data_out_valid(stream_blocks_8_attention_key_weight_valid)
);

stream_blocks_8_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_8_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_8_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_8_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_8_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_attention_mkey_bias),
    .edata_out(stream_blocks_8_attention_ekey_bias),
    .data_out_ready(stream_blocks_8_attention_key_bias_ready),
    .data_out_valid(stream_blocks_8_attention_key_bias_valid)
);

stream_blocks_8_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_8_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_8_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_attention_mvalue_weight),
    .edata_out(stream_blocks_8_attention_evalue_weight),
    .data_out_ready(stream_blocks_8_attention_value_weight_ready),
    .data_out_valid(stream_blocks_8_attention_value_weight_valid)
);

stream_blocks_8_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_8_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_8_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_8_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_8_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_attention_mvalue_bias),
    .edata_out(stream_blocks_8_attention_evalue_bias),
    .data_out_ready(stream_blocks_8_attention_value_bias_ready),
    .data_out_valid(stream_blocks_8_attention_value_bias_valid)
);

stream_blocks_8_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_8_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_8_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_attention_mproj_weight),
    .edata_out(stream_blocks_8_attention_eproj_weight),
    .data_out_ready(stream_blocks_8_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_8_attention_proj_weight_valid)
);

stream_blocks_8_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_8_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_8_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_8_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_8_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_attention_mproj_bias),
    .edata_out(stream_blocks_8_attention_eproj_bias),
    .data_out_ready(stream_blocks_8_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_8_attention_proj_bias_valid)
);

// stream_blocks_8_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_8_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_8_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_8_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_8_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_8_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_8_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_8_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_8_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_8_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_8_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_8_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_8_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_8_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_8_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_8_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_8_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_8_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_8_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_8_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_8_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_8_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_8_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_8_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_8_norm2_mweight),
    .eweight(stream_blocks_8_norm2_eweight),
    .weight_valid(stream_blocks_8_norm2_weight_valid),
    .weight_ready(stream_blocks_8_norm2_weight_ready),
        
    .mbias(stream_blocks_8_norm2_mbias),
    .ebias(stream_blocks_8_norm2_ebias),
    .bias_valid(stream_blocks_8_norm2_bias_valid),
    .bias_ready(stream_blocks_8_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_8_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_8_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_8_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_8_norm2_data_out_0_ready)
);

stream_blocks_8_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_8_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_8_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_8_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_8_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_8_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_8_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_norm2_mweight),
    .edata_out(stream_blocks_8_norm2_eweight),
    .data_out_ready(stream_blocks_8_norm2_weight_ready),
    .data_out_valid(stream_blocks_8_norm2_weight_valid)
);

stream_blocks_8_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_8_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_8_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_8_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_8_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_8_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_8_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_8_norm2_mbias),
    .edata_out(stream_blocks_8_norm2_ebias),
    .data_out_ready(stream_blocks_8_norm2_bias_ready),
    .data_out_valid(stream_blocks_8_norm2_bias_valid)
);

// stream_blocks_8_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_8_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_8_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_8_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_8_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_8_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_8_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_8_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_8_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_8_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_8_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_8_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_8_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_8_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_8_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_8_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_8_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_8_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_8_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_8_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_8_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_8_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_8_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_8_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_8_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_8_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_8_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_8_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_8_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_8_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_8_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_8_add_1_data_out_0_ready)
);

// fork2_18
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_18_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_18_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_18_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_18_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_18_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_18_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_18_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_18_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_18_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_18_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_18_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_18_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_18_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_18_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_18_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_18_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_18_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_18_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_18_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_18_mdata_in_0),
    .edata_in_0(fork2_18_edata_in_0),
    .data_in_0_valid(fork2_18_data_in_0_valid),
    .data_in_0_ready(fork2_18_data_in_0_ready),
        
    .mdata_out_0(fork2_18_mdata_out_0),
    .edata_out_0(fork2_18_edata_out_0),
    .data_out_0_valid(fork2_18_data_out_0_valid),
    .data_out_0_ready(fork2_18_data_out_0_ready),
        
    .mdata_out_1(fork2_18_mdata_out_1),
    .edata_out_1(fork2_18_edata_out_1),
    .data_out_1_valid(fork2_18_data_out_1_valid),
    .data_out_1_ready(fork2_18_data_out_1_ready)
);

// stream_blocks_9_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_9_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_9_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_9_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_9_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_9_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_9_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_9_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_9_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_9_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_9_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_9_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_9_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_9_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_9_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_9_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_9_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_9_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_9_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_9_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_9_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_9_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_9_linear1_mweight),
    .eweight(stream_blocks_9_linear1_eweight),
    .weight_valid(stream_blocks_9_linear1_weight_valid),
    .weight_ready(stream_blocks_9_linear1_weight_ready),
        
    .mbias(stream_blocks_9_linear1_mbias),
    .ebias(stream_blocks_9_linear1_ebias),
    .bias_valid(stream_blocks_9_linear1_bias_valid),
    .bias_ready(stream_blocks_9_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_9_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_9_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_9_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_9_linear1_data_out_0_ready)
);

stream_blocks_9_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_9_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_9_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_9_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_linear1_mweight),
    .edata_out(stream_blocks_9_linear1_eweight),
    .data_out_ready(stream_blocks_9_linear1_weight_ready),
    .data_out_valid(stream_blocks_9_linear1_weight_valid)
);

stream_blocks_9_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_9_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_9_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_9_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_9_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_linear1_mbias),
    .edata_out(stream_blocks_9_linear1_ebias),
    .data_out_ready(stream_blocks_9_linear1_bias_ready),
    .data_out_valid(stream_blocks_9_linear1_bias_valid)
);

// stream_blocks_9_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_9_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_9_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_9_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_9_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_9_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_9_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_9_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_9_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_9_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_9_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_9_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_9_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_9_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_9_act_mdata_in_0),
    .edata_in_0(stream_blocks_9_act_edata_in_0),
    .data_in_0_valid(stream_blocks_9_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_9_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_9_act_mdata_out_0),
    .edata_out_0(stream_blocks_9_act_edata_out_0),
    .data_out_0_valid(stream_blocks_9_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_9_act_data_out_0_ready)
);

// stream_blocks_9_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_9_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_9_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_9_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_9_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_9_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_9_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_9_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_9_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_9_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_9_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_9_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_9_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_9_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_9_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_9_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_9_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_9_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_9_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_9_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_9_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_9_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_9_linear2_mweight),
    .eweight(stream_blocks_9_linear2_eweight),
    .weight_valid(stream_blocks_9_linear2_weight_valid),
    .weight_ready(stream_blocks_9_linear2_weight_ready),
        
    .mbias(stream_blocks_9_linear2_mbias),
    .ebias(stream_blocks_9_linear2_ebias),
    .bias_valid(stream_blocks_9_linear2_bias_valid),
    .bias_ready(stream_blocks_9_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_9_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_9_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_9_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_9_linear2_data_out_0_ready)
);

stream_blocks_9_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_9_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_9_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_9_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_linear2_mweight),
    .edata_out(stream_blocks_9_linear2_eweight),
    .data_out_ready(stream_blocks_9_linear2_weight_ready),
    .data_out_valid(stream_blocks_9_linear2_weight_valid)
);

stream_blocks_9_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_9_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_9_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_9_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_9_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_linear2_mbias),
    .edata_out(stream_blocks_9_linear2_ebias),
    .data_out_ready(stream_blocks_9_linear2_bias_ready),
    .data_out_valid(stream_blocks_9_linear2_bias_valid)
);

// stream_blocks_9_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_9_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_9_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_9_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_9_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_9_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_9_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_9_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_9_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_9_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_9_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_9_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_9_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_9_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_9_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_9_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_9_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_9_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_9_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_9_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_9_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_9_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_9_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_9_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_9_norm1_mweight),
    .eweight(stream_blocks_9_norm1_eweight),
    .weight_valid(stream_blocks_9_norm1_weight_valid),
    .weight_ready(stream_blocks_9_norm1_weight_ready),
        
    .mbias(stream_blocks_9_norm1_mbias),
    .ebias(stream_blocks_9_norm1_ebias),
    .bias_valid(stream_blocks_9_norm1_bias_valid),
    .bias_ready(stream_blocks_9_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_9_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_9_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_9_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_9_norm1_data_out_0_ready)
);

stream_blocks_9_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_9_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_9_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_9_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_norm1_mweight),
    .edata_out(stream_blocks_9_norm1_eweight),
    .data_out_ready(stream_blocks_9_norm1_weight_ready),
    .data_out_valid(stream_blocks_9_norm1_weight_valid)
);

stream_blocks_9_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_9_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_9_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_9_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_9_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_norm1_mbias),
    .edata_out(stream_blocks_9_norm1_ebias),
    .data_out_ready(stream_blocks_9_norm1_bias_ready),
    .data_out_valid(stream_blocks_9_norm1_bias_valid)
);

// stream_blocks_9_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_9_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_9_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_9_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_9_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_9_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_9_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_9_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_9_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_9_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_9_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_9_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_9_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_9_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_9_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_9_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_9_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_9_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_9_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_9_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_9_add_mdata_in_0),
    .edata_in_0(stream_blocks_9_add_edata_in_0),
    .data_in_0_valid(stream_blocks_9_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_9_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_9_add_mdata_in_1),
    .edata_in_1(stream_blocks_9_add_edata_in_1),
    .data_in_1_valid(stream_blocks_9_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_9_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_9_add_mdata_out_0),
    .edata_out_0(stream_blocks_9_add_edata_out_0),
    .data_out_0_valid(stream_blocks_9_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_9_add_data_out_0_ready)
);

// fork2_19
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_19_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_19_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_19_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_19_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_19_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_19_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_19_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_19_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_19_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_19_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_19_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_19_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_19_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_19_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_19_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_19_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_19_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_19_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_19_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_19_mdata_in_0),
    .edata_in_0(fork2_19_edata_in_0),
    .data_in_0_valid(fork2_19_data_in_0_valid),
    .data_in_0_ready(fork2_19_data_in_0_ready),
        
    .mdata_out_0(fork2_19_mdata_out_0),
    .edata_out_0(fork2_19_edata_out_0),
    .data_out_0_valid(fork2_19_data_out_0_valid),
    .data_out_0_ready(fork2_19_data_out_0_ready),
        
    .mdata_out_1(fork2_19_mdata_out_1),
    .edata_out_1(fork2_19_edata_out_1),
    .data_out_1_valid(fork2_19_data_out_1_valid),
    .data_out_1_ready(fork2_19_data_out_1_ready)
);

// stream_blocks_9_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_9_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_9_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_9_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_9_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_9_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_9_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_9_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_9_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_9_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_9_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_9_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_9_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_9_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_9_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_9_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_9_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_9_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_9_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_9_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_9_attention_mdata_in_0),
    .edata_in_0(stream_blocks_9_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_9_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_9_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_9_attention_mquery_weight),
    .equery_weight(stream_blocks_9_attention_equery_weight),
    .query_weight_valid(stream_blocks_9_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_9_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_9_attention_mquery_bias),
    .equery_bias(stream_blocks_9_attention_equery_bias),
    .query_bias_valid(stream_blocks_9_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_9_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_9_attention_mkey_weight),
    .ekey_weight(stream_blocks_9_attention_ekey_weight),
    .key_weight_valid(stream_blocks_9_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_9_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_9_attention_mkey_bias),
    .ekey_bias(stream_blocks_9_attention_ekey_bias),
    .key_bias_valid(stream_blocks_9_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_9_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_9_attention_mvalue_weight),
    .evalue_weight(stream_blocks_9_attention_evalue_weight),
    .value_weight_valid(stream_blocks_9_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_9_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_9_attention_mvalue_bias),
    .evalue_bias(stream_blocks_9_attention_evalue_bias),
    .value_bias_valid(stream_blocks_9_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_9_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_9_attention_mproj_weight),
    .eproj_weight(stream_blocks_9_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_9_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_9_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_9_attention_mproj_bias),
    .eproj_bias(stream_blocks_9_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_9_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_9_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_9_attention_mdata_out_0),
    .edata_out_0(stream_blocks_9_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_9_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_9_attention_data_out_0_ready)
);

stream_blocks_9_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_9_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_9_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_attention_mquery_weight),
    .edata_out(stream_blocks_9_attention_equery_weight),
    .data_out_ready(stream_blocks_9_attention_query_weight_ready),
    .data_out_valid(stream_blocks_9_attention_query_weight_valid)
);

stream_blocks_9_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_9_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_9_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_9_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_9_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_attention_mquery_bias),
    .edata_out(stream_blocks_9_attention_equery_bias),
    .data_out_ready(stream_blocks_9_attention_query_bias_ready),
    .data_out_valid(stream_blocks_9_attention_query_bias_valid)
);

stream_blocks_9_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_9_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_9_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_9_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_attention_mkey_weight),
    .edata_out(stream_blocks_9_attention_ekey_weight),
    .data_out_ready(stream_blocks_9_attention_key_weight_ready),
    .data_out_valid(stream_blocks_9_attention_key_weight_valid)
);

stream_blocks_9_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_9_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_9_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_9_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_9_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_attention_mkey_bias),
    .edata_out(stream_blocks_9_attention_ekey_bias),
    .data_out_ready(stream_blocks_9_attention_key_bias_ready),
    .data_out_valid(stream_blocks_9_attention_key_bias_valid)
);

stream_blocks_9_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_9_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_9_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_attention_mvalue_weight),
    .edata_out(stream_blocks_9_attention_evalue_weight),
    .data_out_ready(stream_blocks_9_attention_value_weight_ready),
    .data_out_valid(stream_blocks_9_attention_value_weight_valid)
);

stream_blocks_9_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_9_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_9_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_9_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_9_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_attention_mvalue_bias),
    .edata_out(stream_blocks_9_attention_evalue_bias),
    .data_out_ready(stream_blocks_9_attention_value_bias_ready),
    .data_out_valid(stream_blocks_9_attention_value_bias_valid)
);

stream_blocks_9_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_9_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_9_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_attention_mproj_weight),
    .edata_out(stream_blocks_9_attention_eproj_weight),
    .data_out_ready(stream_blocks_9_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_9_attention_proj_weight_valid)
);

stream_blocks_9_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_9_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_9_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_9_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_9_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_attention_mproj_bias),
    .edata_out(stream_blocks_9_attention_eproj_bias),
    .data_out_ready(stream_blocks_9_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_9_attention_proj_bias_valid)
);

// stream_blocks_9_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_9_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_9_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_9_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_9_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_9_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_9_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_9_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_9_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_9_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_9_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_9_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_9_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_9_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_9_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_9_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_9_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_9_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_9_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_9_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_9_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_9_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_9_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_9_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_9_norm2_mweight),
    .eweight(stream_blocks_9_norm2_eweight),
    .weight_valid(stream_blocks_9_norm2_weight_valid),
    .weight_ready(stream_blocks_9_norm2_weight_ready),
        
    .mbias(stream_blocks_9_norm2_mbias),
    .ebias(stream_blocks_9_norm2_ebias),
    .bias_valid(stream_blocks_9_norm2_bias_valid),
    .bias_ready(stream_blocks_9_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_9_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_9_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_9_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_9_norm2_data_out_0_ready)
);

stream_blocks_9_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_9_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_9_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_9_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_9_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_9_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_9_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_norm2_mweight),
    .edata_out(stream_blocks_9_norm2_eweight),
    .data_out_ready(stream_blocks_9_norm2_weight_ready),
    .data_out_valid(stream_blocks_9_norm2_weight_valid)
);

stream_blocks_9_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_9_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_9_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_9_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_9_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_9_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_9_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_9_norm2_mbias),
    .edata_out(stream_blocks_9_norm2_ebias),
    .data_out_ready(stream_blocks_9_norm2_bias_ready),
    .data_out_valid(stream_blocks_9_norm2_bias_valid)
);

// stream_blocks_9_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_9_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_9_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_9_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_9_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_9_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_9_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_9_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_9_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_9_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_9_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_9_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_9_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_9_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_9_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_9_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_9_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_9_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_9_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_9_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_9_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_9_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_9_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_9_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_9_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_9_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_9_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_9_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_9_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_9_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_9_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_9_add_1_data_out_0_ready)
);

// fork2_20
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_20_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_20_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_20_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_20_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_20_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_20_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_20_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_20_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_20_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_20_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_20_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_20_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_20_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_20_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_20_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_20_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_20_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_20_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_20_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_20_mdata_in_0),
    .edata_in_0(fork2_20_edata_in_0),
    .data_in_0_valid(fork2_20_data_in_0_valid),
    .data_in_0_ready(fork2_20_data_in_0_ready),
        
    .mdata_out_0(fork2_20_mdata_out_0),
    .edata_out_0(fork2_20_edata_out_0),
    .data_out_0_valid(fork2_20_data_out_0_valid),
    .data_out_0_ready(fork2_20_data_out_0_ready),
        
    .mdata_out_1(fork2_20_mdata_out_1),
    .edata_out_1(fork2_20_edata_out_1),
    .data_out_1_valid(fork2_20_data_out_1_valid),
    .data_out_1_ready(fork2_20_data_out_1_ready)
);

// stream_blocks_10_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_10_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_10_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_10_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_10_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_10_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_10_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_10_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_10_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_10_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_10_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_10_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_10_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_10_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_10_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_10_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_10_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_10_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_10_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_10_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_10_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_10_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_10_linear1_mweight),
    .eweight(stream_blocks_10_linear1_eweight),
    .weight_valid(stream_blocks_10_linear1_weight_valid),
    .weight_ready(stream_blocks_10_linear1_weight_ready),
        
    .mbias(stream_blocks_10_linear1_mbias),
    .ebias(stream_blocks_10_linear1_ebias),
    .bias_valid(stream_blocks_10_linear1_bias_valid),
    .bias_ready(stream_blocks_10_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_10_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_10_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_10_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_10_linear1_data_out_0_ready)
);

stream_blocks_10_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_10_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_10_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_10_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_linear1_mweight),
    .edata_out(stream_blocks_10_linear1_eweight),
    .data_out_ready(stream_blocks_10_linear1_weight_ready),
    .data_out_valid(stream_blocks_10_linear1_weight_valid)
);

stream_blocks_10_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_10_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_10_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_10_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_10_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_linear1_mbias),
    .edata_out(stream_blocks_10_linear1_ebias),
    .data_out_ready(stream_blocks_10_linear1_bias_ready),
    .data_out_valid(stream_blocks_10_linear1_bias_valid)
);

// stream_blocks_10_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_10_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_10_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_10_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_10_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_10_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_10_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_10_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_10_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_10_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_10_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_10_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_10_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_10_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_10_act_mdata_in_0),
    .edata_in_0(stream_blocks_10_act_edata_in_0),
    .data_in_0_valid(stream_blocks_10_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_10_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_10_act_mdata_out_0),
    .edata_out_0(stream_blocks_10_act_edata_out_0),
    .data_out_0_valid(stream_blocks_10_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_10_act_data_out_0_ready)
);

// stream_blocks_10_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_10_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_10_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_10_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_10_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_10_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_10_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_10_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_10_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_10_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_10_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_10_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_10_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_10_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_10_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_10_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_10_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_10_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_10_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_10_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_10_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_10_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_10_linear2_mweight),
    .eweight(stream_blocks_10_linear2_eweight),
    .weight_valid(stream_blocks_10_linear2_weight_valid),
    .weight_ready(stream_blocks_10_linear2_weight_ready),
        
    .mbias(stream_blocks_10_linear2_mbias),
    .ebias(stream_blocks_10_linear2_ebias),
    .bias_valid(stream_blocks_10_linear2_bias_valid),
    .bias_ready(stream_blocks_10_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_10_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_10_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_10_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_10_linear2_data_out_0_ready)
);

stream_blocks_10_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_10_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_10_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_10_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_linear2_mweight),
    .edata_out(stream_blocks_10_linear2_eweight),
    .data_out_ready(stream_blocks_10_linear2_weight_ready),
    .data_out_valid(stream_blocks_10_linear2_weight_valid)
);

stream_blocks_10_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_10_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_10_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_10_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_10_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_linear2_mbias),
    .edata_out(stream_blocks_10_linear2_ebias),
    .data_out_ready(stream_blocks_10_linear2_bias_ready),
    .data_out_valid(stream_blocks_10_linear2_bias_valid)
);

// stream_blocks_10_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_10_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_10_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_10_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_10_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_10_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_10_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_10_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_10_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_10_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_10_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_10_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_10_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_10_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_10_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_10_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_10_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_10_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_10_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_10_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_10_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_10_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_10_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_10_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_10_norm1_mweight),
    .eweight(stream_blocks_10_norm1_eweight),
    .weight_valid(stream_blocks_10_norm1_weight_valid),
    .weight_ready(stream_blocks_10_norm1_weight_ready),
        
    .mbias(stream_blocks_10_norm1_mbias),
    .ebias(stream_blocks_10_norm1_ebias),
    .bias_valid(stream_blocks_10_norm1_bias_valid),
    .bias_ready(stream_blocks_10_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_10_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_10_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_10_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_10_norm1_data_out_0_ready)
);

stream_blocks_10_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_10_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_10_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_10_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_norm1_mweight),
    .edata_out(stream_blocks_10_norm1_eweight),
    .data_out_ready(stream_blocks_10_norm1_weight_ready),
    .data_out_valid(stream_blocks_10_norm1_weight_valid)
);

stream_blocks_10_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_10_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_10_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_10_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_10_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_norm1_mbias),
    .edata_out(stream_blocks_10_norm1_ebias),
    .data_out_ready(stream_blocks_10_norm1_bias_ready),
    .data_out_valid(stream_blocks_10_norm1_bias_valid)
);

// stream_blocks_10_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_10_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_10_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_10_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_10_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_10_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_10_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_10_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_10_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_10_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_10_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_10_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_10_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_10_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_10_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_10_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_10_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_10_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_10_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_10_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_10_add_mdata_in_0),
    .edata_in_0(stream_blocks_10_add_edata_in_0),
    .data_in_0_valid(stream_blocks_10_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_10_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_10_add_mdata_in_1),
    .edata_in_1(stream_blocks_10_add_edata_in_1),
    .data_in_1_valid(stream_blocks_10_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_10_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_10_add_mdata_out_0),
    .edata_out_0(stream_blocks_10_add_edata_out_0),
    .data_out_0_valid(stream_blocks_10_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_10_add_data_out_0_ready)
);

// fork2_21
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_21_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_21_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_21_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_21_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_21_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_21_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_21_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_21_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_21_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_21_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_21_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_21_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_21_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_21_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_21_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_21_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_21_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_21_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_21_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_21_mdata_in_0),
    .edata_in_0(fork2_21_edata_in_0),
    .data_in_0_valid(fork2_21_data_in_0_valid),
    .data_in_0_ready(fork2_21_data_in_0_ready),
        
    .mdata_out_0(fork2_21_mdata_out_0),
    .edata_out_0(fork2_21_edata_out_0),
    .data_out_0_valid(fork2_21_data_out_0_valid),
    .data_out_0_ready(fork2_21_data_out_0_ready),
        
    .mdata_out_1(fork2_21_mdata_out_1),
    .edata_out_1(fork2_21_edata_out_1),
    .data_out_1_valid(fork2_21_data_out_1_valid),
    .data_out_1_ready(fork2_21_data_out_1_ready)
);

// stream_blocks_10_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_10_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_10_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_10_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_10_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_10_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_10_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_10_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_10_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_10_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_10_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_10_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_10_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_10_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_10_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_10_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_10_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_10_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_10_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_10_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_10_attention_mdata_in_0),
    .edata_in_0(stream_blocks_10_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_10_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_10_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_10_attention_mquery_weight),
    .equery_weight(stream_blocks_10_attention_equery_weight),
    .query_weight_valid(stream_blocks_10_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_10_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_10_attention_mquery_bias),
    .equery_bias(stream_blocks_10_attention_equery_bias),
    .query_bias_valid(stream_blocks_10_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_10_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_10_attention_mkey_weight),
    .ekey_weight(stream_blocks_10_attention_ekey_weight),
    .key_weight_valid(stream_blocks_10_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_10_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_10_attention_mkey_bias),
    .ekey_bias(stream_blocks_10_attention_ekey_bias),
    .key_bias_valid(stream_blocks_10_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_10_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_10_attention_mvalue_weight),
    .evalue_weight(stream_blocks_10_attention_evalue_weight),
    .value_weight_valid(stream_blocks_10_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_10_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_10_attention_mvalue_bias),
    .evalue_bias(stream_blocks_10_attention_evalue_bias),
    .value_bias_valid(stream_blocks_10_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_10_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_10_attention_mproj_weight),
    .eproj_weight(stream_blocks_10_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_10_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_10_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_10_attention_mproj_bias),
    .eproj_bias(stream_blocks_10_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_10_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_10_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_10_attention_mdata_out_0),
    .edata_out_0(stream_blocks_10_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_10_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_10_attention_data_out_0_ready)
);

stream_blocks_10_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_10_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_10_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_attention_mquery_weight),
    .edata_out(stream_blocks_10_attention_equery_weight),
    .data_out_ready(stream_blocks_10_attention_query_weight_ready),
    .data_out_valid(stream_blocks_10_attention_query_weight_valid)
);

stream_blocks_10_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_10_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_10_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_10_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_10_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_attention_mquery_bias),
    .edata_out(stream_blocks_10_attention_equery_bias),
    .data_out_ready(stream_blocks_10_attention_query_bias_ready),
    .data_out_valid(stream_blocks_10_attention_query_bias_valid)
);

stream_blocks_10_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_10_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_10_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_10_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_attention_mkey_weight),
    .edata_out(stream_blocks_10_attention_ekey_weight),
    .data_out_ready(stream_blocks_10_attention_key_weight_ready),
    .data_out_valid(stream_blocks_10_attention_key_weight_valid)
);

stream_blocks_10_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_10_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_10_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_10_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_10_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_attention_mkey_bias),
    .edata_out(stream_blocks_10_attention_ekey_bias),
    .data_out_ready(stream_blocks_10_attention_key_bias_ready),
    .data_out_valid(stream_blocks_10_attention_key_bias_valid)
);

stream_blocks_10_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_10_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_10_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_attention_mvalue_weight),
    .edata_out(stream_blocks_10_attention_evalue_weight),
    .data_out_ready(stream_blocks_10_attention_value_weight_ready),
    .data_out_valid(stream_blocks_10_attention_value_weight_valid)
);

stream_blocks_10_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_10_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_10_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_10_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_10_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_attention_mvalue_bias),
    .edata_out(stream_blocks_10_attention_evalue_bias),
    .data_out_ready(stream_blocks_10_attention_value_bias_ready),
    .data_out_valid(stream_blocks_10_attention_value_bias_valid)
);

stream_blocks_10_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_10_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_10_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_attention_mproj_weight),
    .edata_out(stream_blocks_10_attention_eproj_weight),
    .data_out_ready(stream_blocks_10_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_10_attention_proj_weight_valid)
);

stream_blocks_10_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_10_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_10_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_10_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_10_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_attention_mproj_bias),
    .edata_out(stream_blocks_10_attention_eproj_bias),
    .data_out_ready(stream_blocks_10_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_10_attention_proj_bias_valid)
);

// stream_blocks_10_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_10_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_10_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_10_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_10_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_10_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_10_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_10_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_10_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_10_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_10_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_10_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_10_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_10_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_10_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_10_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_10_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_10_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_10_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_10_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_10_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_10_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_10_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_10_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_10_norm2_mweight),
    .eweight(stream_blocks_10_norm2_eweight),
    .weight_valid(stream_blocks_10_norm2_weight_valid),
    .weight_ready(stream_blocks_10_norm2_weight_ready),
        
    .mbias(stream_blocks_10_norm2_mbias),
    .ebias(stream_blocks_10_norm2_ebias),
    .bias_valid(stream_blocks_10_norm2_bias_valid),
    .bias_ready(stream_blocks_10_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_10_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_10_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_10_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_10_norm2_data_out_0_ready)
);

stream_blocks_10_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_10_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_10_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_10_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_10_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_10_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_10_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_norm2_mweight),
    .edata_out(stream_blocks_10_norm2_eweight),
    .data_out_ready(stream_blocks_10_norm2_weight_ready),
    .data_out_valid(stream_blocks_10_norm2_weight_valid)
);

stream_blocks_10_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_10_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_10_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_10_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_10_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_10_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_10_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_10_norm2_mbias),
    .edata_out(stream_blocks_10_norm2_ebias),
    .data_out_ready(stream_blocks_10_norm2_bias_ready),
    .data_out_valid(stream_blocks_10_norm2_bias_valid)
);

// stream_blocks_10_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_10_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_10_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_10_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_10_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_10_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_10_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_10_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_10_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_10_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_10_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_10_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_10_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_10_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_10_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_10_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_10_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_10_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_10_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_10_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_10_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_10_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_10_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_10_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_10_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_10_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_10_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_10_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_10_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_10_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_10_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_10_add_1_data_out_0_ready)
);

// fork2_22
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_22_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_22_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_22_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_22_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_22_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_22_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_22_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_22_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_22_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_22_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_22_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_22_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_22_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_22_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_22_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_22_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_22_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_22_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_22_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_22_mdata_in_0),
    .edata_in_0(fork2_22_edata_in_0),
    .data_in_0_valid(fork2_22_data_in_0_valid),
    .data_in_0_ready(fork2_22_data_in_0_ready),
        
    .mdata_out_0(fork2_22_mdata_out_0),
    .edata_out_0(fork2_22_edata_out_0),
    .data_out_0_valid(fork2_22_data_out_0_valid),
    .data_out_0_ready(fork2_22_data_out_0_ready),
        
    .mdata_out_1(fork2_22_mdata_out_1),
    .edata_out_1(fork2_22_edata_out_1),
    .data_out_1_valid(fork2_22_data_out_1_valid),
    .data_out_1_ready(fork2_22_data_out_1_ready)
);

// stream_blocks_11_linear1
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_11_linear1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_11_linear1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_11_linear1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_11_linear1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_11_linear1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_11_linear1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_11_linear1_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_11_linear1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_linear1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_linear1_WEIGHT_TENSOR_SIZE_DIM_1), // = 768
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_11_linear1_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_11_linear1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_linear1_BIAS_TENSOR_SIZE_DIM_0), // = 768
    .BIAS_PARALLELISM_DIM_0(stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_linear1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_11_linear1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_11_linear1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_11_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_11_linear1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_11_linear1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_11_linear1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_11_linear1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_11_linear1_mdata_in_0),
    .edata_in_0(stream_blocks_11_linear1_edata_in_0),
    .data_in_0_valid(stream_blocks_11_linear1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_11_linear1_data_in_0_ready),
        
    .mweight(stream_blocks_11_linear1_mweight),
    .eweight(stream_blocks_11_linear1_eweight),
    .weight_valid(stream_blocks_11_linear1_weight_valid),
    .weight_ready(stream_blocks_11_linear1_weight_ready),
        
    .mbias(stream_blocks_11_linear1_mbias),
    .ebias(stream_blocks_11_linear1_ebias),
    .bias_valid(stream_blocks_11_linear1_bias_valid),
    .bias_ready(stream_blocks_11_linear1_bias_ready),
        
    .mdata_out_0(stream_blocks_11_linear1_mdata_out_0),
    .edata_out_0(stream_blocks_11_linear1_edata_out_0),
    .data_out_0_valid(stream_blocks_11_linear1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_11_linear1_data_out_0_ready)
);

stream_blocks_11_linear1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_11_linear1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_11_linear1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_linear1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_linear1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_linear1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_11_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_linear1_mweight),
    .edata_out(stream_blocks_11_linear1_eweight),
    .data_out_ready(stream_blocks_11_linear1_weight_ready),
    .data_out_valid(stream_blocks_11_linear1_weight_valid)
);

stream_blocks_11_linear1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_11_linear1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_11_linear1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_linear1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_linear1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_11_linear1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_11_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_linear1_mbias),
    .edata_out(stream_blocks_11_linear1_ebias),
    .data_out_ready(stream_blocks_11_linear1_bias_ready),
    .data_out_valid(stream_blocks_11_linear1_bias_valid)
);

// stream_blocks_11_act
mxint_gelu #(
    .DATA_IN_0_PRECISION_0(stream_blocks_11_act_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_11_act_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_11_act_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_11_act_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_11_act_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_11_act_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_11_act_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_11_act_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_11_act_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_11_act_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_11_act_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_11_act_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_11_act_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_11_act_mdata_in_0),
    .edata_in_0(stream_blocks_11_act_edata_in_0),
    .data_in_0_valid(stream_blocks_11_act_data_in_0_valid),
    .data_in_0_ready(stream_blocks_11_act_data_in_0_ready),
        
    .mdata_out_0(stream_blocks_11_act_mdata_out_0),
    .edata_out_0(stream_blocks_11_act_edata_out_0),
    .data_out_0_valid(stream_blocks_11_act_data_out_0_valid),
    .data_out_0_ready(stream_blocks_11_act_data_out_0_ready)
);

// stream_blocks_11_linear2
mxint_linear #(
    .DATA_IN_0_PRECISION_0(stream_blocks_11_linear2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_11_linear2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_11_linear2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 768
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_11_linear2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_11_linear2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_11_linear2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_11_linear2_WEIGHT_PRECISION_0), // = 4
    .WEIGHT_PRECISION_1(stream_blocks_11_linear2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_linear2_WEIGHT_TENSOR_SIZE_DIM_0), // = 768
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_linear2_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_1), // = 4
    .BIAS_PRECISION_0(stream_blocks_11_linear2_BIAS_PRECISION_0), // = 4
    .BIAS_PRECISION_1(stream_blocks_11_linear2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_linear2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_linear2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_11_linear2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_11_linear2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_11_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_11_linear2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_11_linear2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_11_linear2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_11_linear2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_11_linear2_mdata_in_0),
    .edata_in_0(stream_blocks_11_linear2_edata_in_0),
    .data_in_0_valid(stream_blocks_11_linear2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_11_linear2_data_in_0_ready),
        
    .mweight(stream_blocks_11_linear2_mweight),
    .eweight(stream_blocks_11_linear2_eweight),
    .weight_valid(stream_blocks_11_linear2_weight_valid),
    .weight_ready(stream_blocks_11_linear2_weight_ready),
        
    .mbias(stream_blocks_11_linear2_mbias),
    .ebias(stream_blocks_11_linear2_ebias),
    .bias_valid(stream_blocks_11_linear2_bias_valid),
    .bias_ready(stream_blocks_11_linear2_bias_ready),
        
    .mdata_out_0(stream_blocks_11_linear2_mdata_out_0),
    .edata_out_0(stream_blocks_11_linear2_edata_out_0),
    .data_out_0_valid(stream_blocks_11_linear2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_11_linear2_data_out_0_ready)
);

stream_blocks_11_linear2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_11_linear2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_11_linear2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_linear2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_linear2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_linear2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_11_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_linear2_mweight),
    .edata_out(stream_blocks_11_linear2_eweight),
    .data_out_ready(stream_blocks_11_linear2_weight_ready),
    .data_out_valid(stream_blocks_11_linear2_weight_valid)
);

stream_blocks_11_linear2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_11_linear2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_11_linear2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_linear2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_linear2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_11_linear2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_11_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_linear2_mbias),
    .edata_out(stream_blocks_11_linear2_ebias),
    .data_out_ready(stream_blocks_11_linear2_bias_ready),
    .data_out_valid(stream_blocks_11_linear2_bias_valid)
);

// stream_blocks_11_norm1
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_11_norm1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_11_norm1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_11_norm1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_11_norm1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_11_norm1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_11_norm1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_11_norm1_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_11_norm1_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_norm1_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_norm1_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_11_norm1_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_11_norm1_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_norm1_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_norm1_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_11_norm1_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_11_norm1_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_11_norm1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_11_norm1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_11_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_11_norm1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_11_norm1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_11_norm1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_11_norm1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_11_norm1_mdata_in_0),
    .edata_in_0(stream_blocks_11_norm1_edata_in_0),
    .data_in_0_valid(stream_blocks_11_norm1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_11_norm1_data_in_0_ready),
        
    .mweight(stream_blocks_11_norm1_mweight),
    .eweight(stream_blocks_11_norm1_eweight),
    .weight_valid(stream_blocks_11_norm1_weight_valid),
    .weight_ready(stream_blocks_11_norm1_weight_ready),
        
    .mbias(stream_blocks_11_norm1_mbias),
    .ebias(stream_blocks_11_norm1_ebias),
    .bias_valid(stream_blocks_11_norm1_bias_valid),
    .bias_ready(stream_blocks_11_norm1_bias_ready),
        
    .mdata_out_0(stream_blocks_11_norm1_mdata_out_0),
    .edata_out_0(stream_blocks_11_norm1_edata_out_0),
    .data_out_0_valid(stream_blocks_11_norm1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_11_norm1_data_out_0_ready)
);

stream_blocks_11_norm1_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_11_norm1_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_11_norm1_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_norm1_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_norm1_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_norm1_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_11_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_norm1_mweight),
    .edata_out(stream_blocks_11_norm1_eweight),
    .data_out_ready(stream_blocks_11_norm1_weight_ready),
    .data_out_valid(stream_blocks_11_norm1_weight_valid)
);

stream_blocks_11_norm1_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_11_norm1_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_11_norm1_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_norm1_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_norm1_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_11_norm1_BIAS_PARALLELISM_DIM_1)
) stream_blocks_11_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_norm1_mbias),
    .edata_out(stream_blocks_11_norm1_ebias),
    .data_out_ready(stream_blocks_11_norm1_bias_ready),
    .data_out_valid(stream_blocks_11_norm1_bias_valid)
);

// stream_blocks_11_add
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_11_add_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_11_add_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_11_add_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_11_add_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_11_add_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_11_add_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_11_add_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_11_add_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_11_add_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_11_add_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_11_add_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_11_add_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_11_add_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_11_add_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_11_add_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_11_add_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_11_add_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_11_add_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_11_add_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_11_add_mdata_in_0),
    .edata_in_0(stream_blocks_11_add_edata_in_0),
    .data_in_0_valid(stream_blocks_11_add_data_in_0_valid),
    .data_in_0_ready(stream_blocks_11_add_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_11_add_mdata_in_1),
    .edata_in_1(stream_blocks_11_add_edata_in_1),
    .data_in_1_valid(stream_blocks_11_add_data_in_1_valid),
    .data_in_1_ready(stream_blocks_11_add_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_11_add_mdata_out_0),
    .edata_out_0(stream_blocks_11_add_edata_out_0),
    .data_out_0_valid(stream_blocks_11_add_data_out_0_valid),
    .data_out_0_ready(stream_blocks_11_add_data_out_0_ready)
);

// fork2_23
mxint_fork2 #(
    .DATA_IN_0_PRECISION_0(fork2_23_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(fork2_23_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(fork2_23_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(fork2_23_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(fork2_23_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(fork2_23_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(fork2_23_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(fork2_23_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(fork2_23_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(fork2_23_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(fork2_23_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(fork2_23_DATA_OUT_0_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_1_PRECISION_0(fork2_23_DATA_OUT_1_PRECISION_0), // = 6
    .DATA_OUT_1_PRECISION_1(fork2_23_DATA_OUT_1_PRECISION_1), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_0(fork2_23_DATA_OUT_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_1_PARALLELISM_DIM_0(fork2_23_DATA_OUT_1_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_1_TENSOR_SIZE_DIM_1(fork2_23_DATA_OUT_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_1_PARALLELISM_DIM_1(fork2_23_DATA_OUT_1_PARALLELISM_DIM_1)
) fork2_23_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(fork2_23_mdata_in_0),
    .edata_in_0(fork2_23_edata_in_0),
    .data_in_0_valid(fork2_23_data_in_0_valid),
    .data_in_0_ready(fork2_23_data_in_0_ready),
        
    .mdata_out_0(fork2_23_mdata_out_0),
    .edata_out_0(fork2_23_edata_out_0),
    .data_out_0_valid(fork2_23_data_out_0_valid),
    .data_out_0_ready(fork2_23_data_out_0_ready),
        
    .mdata_out_1(fork2_23_mdata_out_1),
    .edata_out_1(fork2_23_edata_out_1),
    .data_out_1_valid(fork2_23_data_out_1_valid),
    .data_out_1_ready(fork2_23_data_out_1_ready)
);

// stream_blocks_11_attention
mxint_vit_attention_wrap #(
    .DATA_IN_0_PRECISION_0(stream_blocks_11_attention_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_11_attention_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_11_attention_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_11_attention_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_0), // = 6
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_1), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .QUERY_BIAS_PRECISION_0(stream_blocks_11_attention_QUERY_BIAS_PRECISION_0), // = 6
    .QUERY_BIAS_PRECISION_1(stream_blocks_11_attention_QUERY_BIAS_PRECISION_1), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_0), // = 4
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_1), // = 1
    .KEY_WEIGHT_PRECISION_0(stream_blocks_11_attention_KEY_WEIGHT_PRECISION_0), // = 6
    .KEY_WEIGHT_PRECISION_1(stream_blocks_11_attention_KEY_WEIGHT_PRECISION_1), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_0), // = 4
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_1), // = 4
    .KEY_BIAS_PRECISION_0(stream_blocks_11_attention_KEY_BIAS_PRECISION_0), // = 6
    .KEY_BIAS_PRECISION_1(stream_blocks_11_attention_KEY_BIAS_PRECISION_1), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_KEY_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_0), // = 4
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_KEY_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_1), // = 1
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_0), // = 6
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_1), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_0), // = 4
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_1), // = 4
    .VALUE_BIAS_PRECISION_0(stream_blocks_11_attention_VALUE_BIAS_PRECISION_0), // = 6
    .VALUE_BIAS_PRECISION_1(stream_blocks_11_attention_VALUE_BIAS_PRECISION_1), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_0), // = 4
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_1), // = 1
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_0), // = 6
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_1), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_0), // = 4
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1), // = 192
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_1), // = 4
    .PROJ_BIAS_PRECISION_0(stream_blocks_11_attention_PROJ_BIAS_PRECISION_0), // = 6
    .PROJ_BIAS_PRECISION_1(stream_blocks_11_attention_PROJ_BIAS_PRECISION_1), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_0), // = 4
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_11_attention_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_11_attention_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_11_attention_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_11_attention_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_11_attention_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_11_attention_mdata_in_0),
    .edata_in_0(stream_blocks_11_attention_edata_in_0),
    .data_in_0_valid(stream_blocks_11_attention_data_in_0_valid),
    .data_in_0_ready(stream_blocks_11_attention_data_in_0_ready),
        
    .mquery_weight(stream_blocks_11_attention_mquery_weight),
    .equery_weight(stream_blocks_11_attention_equery_weight),
    .query_weight_valid(stream_blocks_11_attention_query_weight_valid),
    .query_weight_ready(stream_blocks_11_attention_query_weight_ready),
        
    .mquery_bias(stream_blocks_11_attention_mquery_bias),
    .equery_bias(stream_blocks_11_attention_equery_bias),
    .query_bias_valid(stream_blocks_11_attention_query_bias_valid),
    .query_bias_ready(stream_blocks_11_attention_query_bias_ready),
        
    .mkey_weight(stream_blocks_11_attention_mkey_weight),
    .ekey_weight(stream_blocks_11_attention_ekey_weight),
    .key_weight_valid(stream_blocks_11_attention_key_weight_valid),
    .key_weight_ready(stream_blocks_11_attention_key_weight_ready),
        
    .mkey_bias(stream_blocks_11_attention_mkey_bias),
    .ekey_bias(stream_blocks_11_attention_ekey_bias),
    .key_bias_valid(stream_blocks_11_attention_key_bias_valid),
    .key_bias_ready(stream_blocks_11_attention_key_bias_ready),
        
    .mvalue_weight(stream_blocks_11_attention_mvalue_weight),
    .evalue_weight(stream_blocks_11_attention_evalue_weight),
    .value_weight_valid(stream_blocks_11_attention_value_weight_valid),
    .value_weight_ready(stream_blocks_11_attention_value_weight_ready),
        
    .mvalue_bias(stream_blocks_11_attention_mvalue_bias),
    .evalue_bias(stream_blocks_11_attention_evalue_bias),
    .value_bias_valid(stream_blocks_11_attention_value_bias_valid),
    .value_bias_ready(stream_blocks_11_attention_value_bias_ready),
        
    .mproj_weight(stream_blocks_11_attention_mproj_weight),
    .eproj_weight(stream_blocks_11_attention_eproj_weight),
    .proj_weight_valid(stream_blocks_11_attention_proj_weight_valid),
    .proj_weight_ready(stream_blocks_11_attention_proj_weight_ready),
        
    .mproj_bias(stream_blocks_11_attention_mproj_bias),
    .eproj_bias(stream_blocks_11_attention_eproj_bias),
    .proj_bias_valid(stream_blocks_11_attention_proj_bias_valid),
    .proj_bias_ready(stream_blocks_11_attention_proj_bias_ready),
        
    .mdata_out_0(stream_blocks_11_attention_mdata_out_0),
    .edata_out_0(stream_blocks_11_attention_edata_out_0),
    .data_out_0_valid(stream_blocks_11_attention_data_out_0_valid),
    .data_out_0_ready(stream_blocks_11_attention_data_out_0_ready)
);

stream_blocks_11_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(stream_blocks_11_attention_QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_attention_QUERY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_11_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_attention_mquery_weight),
    .edata_out(stream_blocks_11_attention_equery_weight),
    .data_out_ready(stream_blocks_11_attention_query_weight_ready),
    .data_out_valid(stream_blocks_11_attention_query_weight_valid)
);

stream_blocks_11_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(stream_blocks_11_attention_QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(stream_blocks_11_attention_QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(stream_blocks_11_attention_QUERY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_11_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_attention_mquery_bias),
    .edata_out(stream_blocks_11_attention_equery_bias),
    .data_out_ready(stream_blocks_11_attention_query_bias_ready),
    .data_out_valid(stream_blocks_11_attention_query_bias_valid)
);

stream_blocks_11_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(stream_blocks_11_attention_KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(stream_blocks_11_attention_KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_attention_KEY_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_11_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_attention_mkey_weight),
    .edata_out(stream_blocks_11_attention_ekey_weight),
    .data_out_ready(stream_blocks_11_attention_key_weight_ready),
    .data_out_valid(stream_blocks_11_attention_key_weight_valid)
);

stream_blocks_11_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(stream_blocks_11_attention_KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(stream_blocks_11_attention_KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(stream_blocks_11_attention_KEY_BIAS_PARALLELISM_DIM_1)
) stream_blocks_11_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_attention_mkey_bias),
    .edata_out(stream_blocks_11_attention_ekey_bias),
    .data_out_ready(stream_blocks_11_attention_key_bias_ready),
    .data_out_valid(stream_blocks_11_attention_key_bias_valid)
);

stream_blocks_11_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(stream_blocks_11_attention_VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_attention_VALUE_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_11_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_attention_mvalue_weight),
    .edata_out(stream_blocks_11_attention_evalue_weight),
    .data_out_ready(stream_blocks_11_attention_value_weight_ready),
    .data_out_valid(stream_blocks_11_attention_value_weight_valid)
);

stream_blocks_11_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(stream_blocks_11_attention_VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(stream_blocks_11_attention_VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(stream_blocks_11_attention_VALUE_BIAS_PARALLELISM_DIM_1)
) stream_blocks_11_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_attention_mvalue_bias),
    .edata_out(stream_blocks_11_attention_evalue_bias),
    .data_out_ready(stream_blocks_11_attention_value_bias_ready),
    .data_out_valid(stream_blocks_11_attention_value_bias_valid)
);

stream_blocks_11_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(stream_blocks_11_attention_PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_attention_PROJ_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_11_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_attention_mproj_weight),
    .edata_out(stream_blocks_11_attention_eproj_weight),
    .data_out_ready(stream_blocks_11_attention_proj_weight_ready),
    .data_out_valid(stream_blocks_11_attention_proj_weight_valid)
);

stream_blocks_11_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(stream_blocks_11_attention_PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(stream_blocks_11_attention_PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_attention_PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_attention_PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(stream_blocks_11_attention_PROJ_BIAS_PARALLELISM_DIM_1)
) stream_blocks_11_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_attention_mproj_bias),
    .edata_out(stream_blocks_11_attention_eproj_bias),
    .data_out_ready(stream_blocks_11_attention_proj_bias_ready),
    .data_out_valid(stream_blocks_11_attention_proj_bias_valid)
);

// stream_blocks_11_norm2
mxint_layernorm #(
    .DATA_IN_0_PRECISION_0(stream_blocks_11_norm2_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_11_norm2_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_11_norm2_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_11_norm2_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_11_norm2_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_11_norm2_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .WEIGHT_PRECISION_0(stream_blocks_11_norm2_WEIGHT_PRECISION_0), // = 6
    .WEIGHT_PRECISION_1(stream_blocks_11_norm2_WEIGHT_PRECISION_1), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_norm2_WEIGHT_TENSOR_SIZE_DIM_0), // = 192
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_0), // = 4
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_norm2_WEIGHT_TENSOR_SIZE_DIM_1), // = 1
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_1), // = 1
    .BIAS_PRECISION_0(stream_blocks_11_norm2_BIAS_PRECISION_0), // = 6
    .BIAS_PRECISION_1(stream_blocks_11_norm2_BIAS_PRECISION_1), // = 4
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_norm2_BIAS_TENSOR_SIZE_DIM_0), // = 192
    .BIAS_PARALLELISM_DIM_0(stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_0), // = 4
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_norm2_BIAS_TENSOR_SIZE_DIM_1), // = 1
    .BIAS_PARALLELISM_DIM_1(stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_1), // = 1
    .ELEMENTWISE_AFFINE(stream_blocks_11_norm2_ELEMENTWISE_AFFINE), // = 1
    .HAS_BIAS(stream_blocks_11_norm2_HAS_BIAS), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_11_norm2_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_11_norm2_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_11_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_11_norm2_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_11_norm2_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_11_norm2_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_11_norm2_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_11_norm2_mdata_in_0),
    .edata_in_0(stream_blocks_11_norm2_edata_in_0),
    .data_in_0_valid(stream_blocks_11_norm2_data_in_0_valid),
    .data_in_0_ready(stream_blocks_11_norm2_data_in_0_ready),
        
    .mweight(stream_blocks_11_norm2_mweight),
    .eweight(stream_blocks_11_norm2_eweight),
    .weight_valid(stream_blocks_11_norm2_weight_valid),
    .weight_ready(stream_blocks_11_norm2_weight_ready),
        
    .mbias(stream_blocks_11_norm2_mbias),
    .ebias(stream_blocks_11_norm2_ebias),
    .bias_valid(stream_blocks_11_norm2_bias_valid),
    .bias_ready(stream_blocks_11_norm2_bias_ready),
        
    .mdata_out_0(stream_blocks_11_norm2_mdata_out_0),
    .edata_out_0(stream_blocks_11_norm2_edata_out_0),
    .data_out_0_valid(stream_blocks_11_norm2_data_out_0_valid),
    .data_out_0_ready(stream_blocks_11_norm2_data_out_0_ready)
);

stream_blocks_11_norm2_weight_source #(
    .WEIGHT_PRECISION_0(stream_blocks_11_norm2_WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(stream_blocks_11_norm2_WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(stream_blocks_11_norm2_WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(stream_blocks_11_norm2_WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(stream_blocks_11_norm2_WEIGHT_PARALLELISM_DIM_1)
) stream_blocks_11_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_norm2_mweight),
    .edata_out(stream_blocks_11_norm2_eweight),
    .data_out_ready(stream_blocks_11_norm2_weight_ready),
    .data_out_valid(stream_blocks_11_norm2_weight_valid)
);

stream_blocks_11_norm2_bias_source #(
    .BIAS_PRECISION_0(stream_blocks_11_norm2_BIAS_PRECISION_0),
    .BIAS_PRECISION_1(stream_blocks_11_norm2_BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(stream_blocks_11_norm2_BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(stream_blocks_11_norm2_BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(stream_blocks_11_norm2_BIAS_PARALLELISM_DIM_1)
) stream_blocks_11_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(stream_blocks_11_norm2_mbias),
    .edata_out(stream_blocks_11_norm2_ebias),
    .data_out_ready(stream_blocks_11_norm2_bias_ready),
    .data_out_valid(stream_blocks_11_norm2_bias_valid)
);

// stream_blocks_11_add_1
mxint_addition #(
    .DATA_IN_0_PRECISION_0(stream_blocks_11_add_1_DATA_IN_0_PRECISION_0), // = 6
    .DATA_IN_0_PRECISION_1(stream_blocks_11_add_1_DATA_IN_0_PRECISION_1), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_0(stream_blocks_11_add_1_DATA_IN_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_0_PARALLELISM_DIM_0(stream_blocks_11_add_1_DATA_IN_0_PARALLELISM_DIM_0), // = 4
    .DATA_IN_0_TENSOR_SIZE_DIM_1(stream_blocks_11_add_1_DATA_IN_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_0_PARALLELISM_DIM_1(stream_blocks_11_add_1_DATA_IN_0_PARALLELISM_DIM_1), // = 1
    .DATA_IN_1_PRECISION_0(stream_blocks_11_add_1_DATA_IN_1_PRECISION_0), // = 6
    .DATA_IN_1_PRECISION_1(stream_blocks_11_add_1_DATA_IN_1_PRECISION_1), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_0(stream_blocks_11_add_1_DATA_IN_1_TENSOR_SIZE_DIM_0), // = 192
    .DATA_IN_1_PARALLELISM_DIM_0(stream_blocks_11_add_1_DATA_IN_1_PARALLELISM_DIM_0), // = 4
    .DATA_IN_1_TENSOR_SIZE_DIM_1(stream_blocks_11_add_1_DATA_IN_1_TENSOR_SIZE_DIM_1), // = 196
    .DATA_IN_1_PARALLELISM_DIM_1(stream_blocks_11_add_1_DATA_IN_1_PARALLELISM_DIM_1), // = 1
    .DATA_OUT_0_PRECISION_0(stream_blocks_11_add_1_DATA_OUT_0_PRECISION_0), // = 6
    .DATA_OUT_0_PRECISION_1(stream_blocks_11_add_1_DATA_OUT_0_PRECISION_1), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_0(stream_blocks_11_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_0), // = 192
    .DATA_OUT_0_PARALLELISM_DIM_0(stream_blocks_11_add_1_DATA_OUT_0_PARALLELISM_DIM_0), // = 4
    .DATA_OUT_0_TENSOR_SIZE_DIM_1(stream_blocks_11_add_1_DATA_OUT_0_TENSOR_SIZE_DIM_1), // = 196
    .DATA_OUT_0_PARALLELISM_DIM_1(stream_blocks_11_add_1_DATA_OUT_0_PARALLELISM_DIM_1)
) stream_blocks_11_add_1_inst (
    .clk(clk),
    .rst(rst),

    .mdata_in_0(stream_blocks_11_add_1_mdata_in_0),
    .edata_in_0(stream_blocks_11_add_1_edata_in_0),
    .data_in_0_valid(stream_blocks_11_add_1_data_in_0_valid),
    .data_in_0_ready(stream_blocks_11_add_1_data_in_0_ready),
        
    .mdata_in_1(stream_blocks_11_add_1_mdata_in_1),
    .edata_in_1(stream_blocks_11_add_1_edata_in_1),
    .data_in_1_valid(stream_blocks_11_add_1_data_in_1_valid),
    .data_in_1_ready(stream_blocks_11_add_1_data_in_1_ready),
        
    .mdata_out_0(stream_blocks_11_add_1_mdata_out_0),
    .edata_out_0(stream_blocks_11_add_1_edata_out_0),
    .data_out_0_valid(stream_blocks_11_add_1_data_out_0_valid),
    .data_out_0_ready(stream_blocks_11_add_1_data_out_0_ready)
);


// --------------------------
//   Interconnections
// --------------------------
    
assign data_in_0_ready = fork2_data_in_0_ready;
assign fork2_data_in_0_valid    = data_in_0_valid;
assign fork2_mdata_in_0    = mdata_in_0;
assign fork2_edata_in_0    = edata_in_0;

assign data_out_0_valid = stream_blocks_11_add_1_data_out_0_valid;
assign stream_blocks_11_add_1_data_out_0_ready    = data_out_0_ready;
assign mdata_out_0 = stream_blocks_11_add_1_mdata_out_0;
assign edata_out_0 = stream_blocks_11_add_1_edata_out_0;

assign fork2_data_out_0_ready  = stream_blocks_0_linear1_data_in_0_ready;
assign stream_blocks_0_linear1_data_in_0_valid    = fork2_data_out_0_valid;
assign stream_blocks_0_linear1_mdata_in_0 = fork2_mdata_out_0;
assign stream_blocks_0_linear1_edata_in_0 = fork2_edata_out_0;

assign stream_blocks_0_linear1_data_out_0_ready  = stream_blocks_0_act_data_in_0_ready;
assign stream_blocks_0_act_data_in_0_valid    = stream_blocks_0_linear1_data_out_0_valid;
assign stream_blocks_0_act_mdata_in_0 = stream_blocks_0_linear1_mdata_out_0;
assign stream_blocks_0_act_edata_in_0 = stream_blocks_0_linear1_edata_out_0;

assign stream_blocks_0_act_data_out_0_ready  = stream_blocks_0_linear2_data_in_0_ready;
assign stream_blocks_0_linear2_data_in_0_valid    = stream_blocks_0_act_data_out_0_valid;
assign stream_blocks_0_linear2_mdata_in_0 = stream_blocks_0_act_mdata_out_0;
assign stream_blocks_0_linear2_edata_in_0 = stream_blocks_0_act_edata_out_0;

assign stream_blocks_0_linear2_data_out_0_ready  = stream_blocks_0_norm1_data_in_0_ready;
assign stream_blocks_0_norm1_data_in_0_valid    = stream_blocks_0_linear2_data_out_0_valid;
assign stream_blocks_0_norm1_mdata_in_0 = stream_blocks_0_linear2_mdata_out_0;
assign stream_blocks_0_norm1_edata_in_0 = stream_blocks_0_linear2_edata_out_0;

assign stream_blocks_0_norm1_data_out_0_ready  = stream_blocks_0_add_data_in_0_ready;
assign stream_blocks_0_add_data_in_0_valid    = stream_blocks_0_norm1_data_out_0_valid;
assign stream_blocks_0_add_mdata_in_0 = stream_blocks_0_norm1_mdata_out_0;
assign stream_blocks_0_add_edata_in_0 = stream_blocks_0_norm1_edata_out_0;

assign fork2_data_out_1_ready  = stream_blocks_0_add_data_in_1_ready;
assign stream_blocks_0_add_data_in_1_valid    = fork2_data_out_1_valid;
assign stream_blocks_0_add_mdata_in_1 = fork2_mdata_out_1;
assign stream_blocks_0_add_edata_in_1 = fork2_edata_out_1;

assign stream_blocks_0_add_data_out_0_ready  = fork2_1_data_in_0_ready;
assign fork2_1_data_in_0_valid    = stream_blocks_0_add_data_out_0_valid;
assign fork2_1_mdata_in_0 = stream_blocks_0_add_mdata_out_0;
assign fork2_1_edata_in_0 = stream_blocks_0_add_edata_out_0;

assign fork2_1_data_out_0_ready  = stream_blocks_0_attention_data_in_0_ready;
assign stream_blocks_0_attention_data_in_0_valid    = fork2_1_data_out_0_valid;
assign stream_blocks_0_attention_mdata_in_0 = fork2_1_mdata_out_0;
assign stream_blocks_0_attention_edata_in_0 = fork2_1_edata_out_0;

assign stream_blocks_0_attention_data_out_0_ready  = stream_blocks_0_norm2_data_in_0_ready;
assign stream_blocks_0_norm2_data_in_0_valid    = stream_blocks_0_attention_data_out_0_valid;
assign stream_blocks_0_norm2_mdata_in_0 = stream_blocks_0_attention_mdata_out_0;
assign stream_blocks_0_norm2_edata_in_0 = stream_blocks_0_attention_edata_out_0;

assign stream_blocks_0_norm2_data_out_0_ready  = stream_blocks_0_add_1_data_in_0_ready;
assign stream_blocks_0_add_1_data_in_0_valid    = stream_blocks_0_norm2_data_out_0_valid;
assign stream_blocks_0_add_1_mdata_in_0 = stream_blocks_0_norm2_mdata_out_0;
assign stream_blocks_0_add_1_edata_in_0 = stream_blocks_0_norm2_edata_out_0;

assign fork2_1_data_out_1_ready  = stream_blocks_0_add_1_data_in_1_ready;
assign stream_blocks_0_add_1_data_in_1_valid    = fork2_1_data_out_1_valid;
assign stream_blocks_0_add_1_mdata_in_1 = fork2_1_mdata_out_1;
assign stream_blocks_0_add_1_edata_in_1 = fork2_1_edata_out_1;

assign stream_blocks_0_add_1_data_out_0_ready  = fork2_2_data_in_0_ready;
assign fork2_2_data_in_0_valid    = stream_blocks_0_add_1_data_out_0_valid;
assign fork2_2_mdata_in_0 = stream_blocks_0_add_1_mdata_out_0;
assign fork2_2_edata_in_0 = stream_blocks_0_add_1_edata_out_0;

assign fork2_2_data_out_0_ready  = stream_blocks_1_linear1_data_in_0_ready;
assign stream_blocks_1_linear1_data_in_0_valid    = fork2_2_data_out_0_valid;
assign stream_blocks_1_linear1_mdata_in_0 = fork2_2_mdata_out_0;
assign stream_blocks_1_linear1_edata_in_0 = fork2_2_edata_out_0;

assign stream_blocks_1_linear1_data_out_0_ready  = stream_blocks_1_act_data_in_0_ready;
assign stream_blocks_1_act_data_in_0_valid    = stream_blocks_1_linear1_data_out_0_valid;
assign stream_blocks_1_act_mdata_in_0 = stream_blocks_1_linear1_mdata_out_0;
assign stream_blocks_1_act_edata_in_0 = stream_blocks_1_linear1_edata_out_0;

assign stream_blocks_1_act_data_out_0_ready  = stream_blocks_1_linear2_data_in_0_ready;
assign stream_blocks_1_linear2_data_in_0_valid    = stream_blocks_1_act_data_out_0_valid;
assign stream_blocks_1_linear2_mdata_in_0 = stream_blocks_1_act_mdata_out_0;
assign stream_blocks_1_linear2_edata_in_0 = stream_blocks_1_act_edata_out_0;

assign stream_blocks_1_linear2_data_out_0_ready  = stream_blocks_1_norm1_data_in_0_ready;
assign stream_blocks_1_norm1_data_in_0_valid    = stream_blocks_1_linear2_data_out_0_valid;
assign stream_blocks_1_norm1_mdata_in_0 = stream_blocks_1_linear2_mdata_out_0;
assign stream_blocks_1_norm1_edata_in_0 = stream_blocks_1_linear2_edata_out_0;

assign stream_blocks_1_norm1_data_out_0_ready  = stream_blocks_1_add_data_in_0_ready;
assign stream_blocks_1_add_data_in_0_valid    = stream_blocks_1_norm1_data_out_0_valid;
assign stream_blocks_1_add_mdata_in_0 = stream_blocks_1_norm1_mdata_out_0;
assign stream_blocks_1_add_edata_in_0 = stream_blocks_1_norm1_edata_out_0;

assign fork2_2_data_out_1_ready  = stream_blocks_1_add_data_in_1_ready;
assign stream_blocks_1_add_data_in_1_valid    = fork2_2_data_out_1_valid;
assign stream_blocks_1_add_mdata_in_1 = fork2_2_mdata_out_1;
assign stream_blocks_1_add_edata_in_1 = fork2_2_edata_out_1;

assign stream_blocks_1_add_data_out_0_ready  = fork2_3_data_in_0_ready;
assign fork2_3_data_in_0_valid    = stream_blocks_1_add_data_out_0_valid;
assign fork2_3_mdata_in_0 = stream_blocks_1_add_mdata_out_0;
assign fork2_3_edata_in_0 = stream_blocks_1_add_edata_out_0;

assign fork2_3_data_out_0_ready  = stream_blocks_1_attention_data_in_0_ready;
assign stream_blocks_1_attention_data_in_0_valid    = fork2_3_data_out_0_valid;
assign stream_blocks_1_attention_mdata_in_0 = fork2_3_mdata_out_0;
assign stream_blocks_1_attention_edata_in_0 = fork2_3_edata_out_0;

assign stream_blocks_1_attention_data_out_0_ready  = stream_blocks_1_norm2_data_in_0_ready;
assign stream_blocks_1_norm2_data_in_0_valid    = stream_blocks_1_attention_data_out_0_valid;
assign stream_blocks_1_norm2_mdata_in_0 = stream_blocks_1_attention_mdata_out_0;
assign stream_blocks_1_norm2_edata_in_0 = stream_blocks_1_attention_edata_out_0;

assign stream_blocks_1_norm2_data_out_0_ready  = stream_blocks_1_add_1_data_in_0_ready;
assign stream_blocks_1_add_1_data_in_0_valid    = stream_blocks_1_norm2_data_out_0_valid;
assign stream_blocks_1_add_1_mdata_in_0 = stream_blocks_1_norm2_mdata_out_0;
assign stream_blocks_1_add_1_edata_in_0 = stream_blocks_1_norm2_edata_out_0;

assign fork2_3_data_out_1_ready  = stream_blocks_1_add_1_data_in_1_ready;
assign stream_blocks_1_add_1_data_in_1_valid    = fork2_3_data_out_1_valid;
assign stream_blocks_1_add_1_mdata_in_1 = fork2_3_mdata_out_1;
assign stream_blocks_1_add_1_edata_in_1 = fork2_3_edata_out_1;

assign stream_blocks_1_add_1_data_out_0_ready  = fork2_4_data_in_0_ready;
assign fork2_4_data_in_0_valid    = stream_blocks_1_add_1_data_out_0_valid;
assign fork2_4_mdata_in_0 = stream_blocks_1_add_1_mdata_out_0;
assign fork2_4_edata_in_0 = stream_blocks_1_add_1_edata_out_0;

assign fork2_4_data_out_0_ready  = stream_blocks_2_linear1_data_in_0_ready;
assign stream_blocks_2_linear1_data_in_0_valid    = fork2_4_data_out_0_valid;
assign stream_blocks_2_linear1_mdata_in_0 = fork2_4_mdata_out_0;
assign stream_blocks_2_linear1_edata_in_0 = fork2_4_edata_out_0;

assign stream_blocks_2_linear1_data_out_0_ready  = stream_blocks_2_act_data_in_0_ready;
assign stream_blocks_2_act_data_in_0_valid    = stream_blocks_2_linear1_data_out_0_valid;
assign stream_blocks_2_act_mdata_in_0 = stream_blocks_2_linear1_mdata_out_0;
assign stream_blocks_2_act_edata_in_0 = stream_blocks_2_linear1_edata_out_0;

assign stream_blocks_2_act_data_out_0_ready  = stream_blocks_2_linear2_data_in_0_ready;
assign stream_blocks_2_linear2_data_in_0_valid    = stream_blocks_2_act_data_out_0_valid;
assign stream_blocks_2_linear2_mdata_in_0 = stream_blocks_2_act_mdata_out_0;
assign stream_blocks_2_linear2_edata_in_0 = stream_blocks_2_act_edata_out_0;

assign stream_blocks_2_linear2_data_out_0_ready  = stream_blocks_2_norm1_data_in_0_ready;
assign stream_blocks_2_norm1_data_in_0_valid    = stream_blocks_2_linear2_data_out_0_valid;
assign stream_blocks_2_norm1_mdata_in_0 = stream_blocks_2_linear2_mdata_out_0;
assign stream_blocks_2_norm1_edata_in_0 = stream_blocks_2_linear2_edata_out_0;

assign stream_blocks_2_norm1_data_out_0_ready  = stream_blocks_2_add_data_in_0_ready;
assign stream_blocks_2_add_data_in_0_valid    = stream_blocks_2_norm1_data_out_0_valid;
assign stream_blocks_2_add_mdata_in_0 = stream_blocks_2_norm1_mdata_out_0;
assign stream_blocks_2_add_edata_in_0 = stream_blocks_2_norm1_edata_out_0;

assign fork2_4_data_out_1_ready  = stream_blocks_2_add_data_in_1_ready;
assign stream_blocks_2_add_data_in_1_valid    = fork2_4_data_out_1_valid;
assign stream_blocks_2_add_mdata_in_1 = fork2_4_mdata_out_1;
assign stream_blocks_2_add_edata_in_1 = fork2_4_edata_out_1;

assign stream_blocks_2_add_data_out_0_ready  = fork2_5_data_in_0_ready;
assign fork2_5_data_in_0_valid    = stream_blocks_2_add_data_out_0_valid;
assign fork2_5_mdata_in_0 = stream_blocks_2_add_mdata_out_0;
assign fork2_5_edata_in_0 = stream_blocks_2_add_edata_out_0;

assign fork2_5_data_out_0_ready  = stream_blocks_2_attention_data_in_0_ready;
assign stream_blocks_2_attention_data_in_0_valid    = fork2_5_data_out_0_valid;
assign stream_blocks_2_attention_mdata_in_0 = fork2_5_mdata_out_0;
assign stream_blocks_2_attention_edata_in_0 = fork2_5_edata_out_0;

assign stream_blocks_2_attention_data_out_0_ready  = stream_blocks_2_norm2_data_in_0_ready;
assign stream_blocks_2_norm2_data_in_0_valid    = stream_blocks_2_attention_data_out_0_valid;
assign stream_blocks_2_norm2_mdata_in_0 = stream_blocks_2_attention_mdata_out_0;
assign stream_blocks_2_norm2_edata_in_0 = stream_blocks_2_attention_edata_out_0;

assign stream_blocks_2_norm2_data_out_0_ready  = stream_blocks_2_add_1_data_in_0_ready;
assign stream_blocks_2_add_1_data_in_0_valid    = stream_blocks_2_norm2_data_out_0_valid;
assign stream_blocks_2_add_1_mdata_in_0 = stream_blocks_2_norm2_mdata_out_0;
assign stream_blocks_2_add_1_edata_in_0 = stream_blocks_2_norm2_edata_out_0;

assign fork2_5_data_out_1_ready  = stream_blocks_2_add_1_data_in_1_ready;
assign stream_blocks_2_add_1_data_in_1_valid    = fork2_5_data_out_1_valid;
assign stream_blocks_2_add_1_mdata_in_1 = fork2_5_mdata_out_1;
assign stream_blocks_2_add_1_edata_in_1 = fork2_5_edata_out_1;

assign stream_blocks_2_add_1_data_out_0_ready  = fork2_6_data_in_0_ready;
assign fork2_6_data_in_0_valid    = stream_blocks_2_add_1_data_out_0_valid;
assign fork2_6_mdata_in_0 = stream_blocks_2_add_1_mdata_out_0;
assign fork2_6_edata_in_0 = stream_blocks_2_add_1_edata_out_0;

assign fork2_6_data_out_0_ready  = stream_blocks_3_linear1_data_in_0_ready;
assign stream_blocks_3_linear1_data_in_0_valid    = fork2_6_data_out_0_valid;
assign stream_blocks_3_linear1_mdata_in_0 = fork2_6_mdata_out_0;
assign stream_blocks_3_linear1_edata_in_0 = fork2_6_edata_out_0;

assign stream_blocks_3_linear1_data_out_0_ready  = stream_blocks_3_act_data_in_0_ready;
assign stream_blocks_3_act_data_in_0_valid    = stream_blocks_3_linear1_data_out_0_valid;
assign stream_blocks_3_act_mdata_in_0 = stream_blocks_3_linear1_mdata_out_0;
assign stream_blocks_3_act_edata_in_0 = stream_blocks_3_linear1_edata_out_0;

assign stream_blocks_3_act_data_out_0_ready  = stream_blocks_3_linear2_data_in_0_ready;
assign stream_blocks_3_linear2_data_in_0_valid    = stream_blocks_3_act_data_out_0_valid;
assign stream_blocks_3_linear2_mdata_in_0 = stream_blocks_3_act_mdata_out_0;
assign stream_blocks_3_linear2_edata_in_0 = stream_blocks_3_act_edata_out_0;

assign stream_blocks_3_linear2_data_out_0_ready  = stream_blocks_3_norm1_data_in_0_ready;
assign stream_blocks_3_norm1_data_in_0_valid    = stream_blocks_3_linear2_data_out_0_valid;
assign stream_blocks_3_norm1_mdata_in_0 = stream_blocks_3_linear2_mdata_out_0;
assign stream_blocks_3_norm1_edata_in_0 = stream_blocks_3_linear2_edata_out_0;

assign stream_blocks_3_norm1_data_out_0_ready  = stream_blocks_3_add_data_in_0_ready;
assign stream_blocks_3_add_data_in_0_valid    = stream_blocks_3_norm1_data_out_0_valid;
assign stream_blocks_3_add_mdata_in_0 = stream_blocks_3_norm1_mdata_out_0;
assign stream_blocks_3_add_edata_in_0 = stream_blocks_3_norm1_edata_out_0;

assign fork2_6_data_out_1_ready  = stream_blocks_3_add_data_in_1_ready;
assign stream_blocks_3_add_data_in_1_valid    = fork2_6_data_out_1_valid;
assign stream_blocks_3_add_mdata_in_1 = fork2_6_mdata_out_1;
assign stream_blocks_3_add_edata_in_1 = fork2_6_edata_out_1;

assign stream_blocks_3_add_data_out_0_ready  = fork2_7_data_in_0_ready;
assign fork2_7_data_in_0_valid    = stream_blocks_3_add_data_out_0_valid;
assign fork2_7_mdata_in_0 = stream_blocks_3_add_mdata_out_0;
assign fork2_7_edata_in_0 = stream_blocks_3_add_edata_out_0;

assign fork2_7_data_out_0_ready  = stream_blocks_3_attention_data_in_0_ready;
assign stream_blocks_3_attention_data_in_0_valid    = fork2_7_data_out_0_valid;
assign stream_blocks_3_attention_mdata_in_0 = fork2_7_mdata_out_0;
assign stream_blocks_3_attention_edata_in_0 = fork2_7_edata_out_0;

assign stream_blocks_3_attention_data_out_0_ready  = stream_blocks_3_norm2_data_in_0_ready;
assign stream_blocks_3_norm2_data_in_0_valid    = stream_blocks_3_attention_data_out_0_valid;
assign stream_blocks_3_norm2_mdata_in_0 = stream_blocks_3_attention_mdata_out_0;
assign stream_blocks_3_norm2_edata_in_0 = stream_blocks_3_attention_edata_out_0;

assign stream_blocks_3_norm2_data_out_0_ready  = stream_blocks_3_add_1_data_in_0_ready;
assign stream_blocks_3_add_1_data_in_0_valid    = stream_blocks_3_norm2_data_out_0_valid;
assign stream_blocks_3_add_1_mdata_in_0 = stream_blocks_3_norm2_mdata_out_0;
assign stream_blocks_3_add_1_edata_in_0 = stream_blocks_3_norm2_edata_out_0;

assign fork2_7_data_out_1_ready  = stream_blocks_3_add_1_data_in_1_ready;
assign stream_blocks_3_add_1_data_in_1_valid    = fork2_7_data_out_1_valid;
assign stream_blocks_3_add_1_mdata_in_1 = fork2_7_mdata_out_1;
assign stream_blocks_3_add_1_edata_in_1 = fork2_7_edata_out_1;

assign stream_blocks_3_add_1_data_out_0_ready  = fork2_8_data_in_0_ready;
assign fork2_8_data_in_0_valid    = stream_blocks_3_add_1_data_out_0_valid;
assign fork2_8_mdata_in_0 = stream_blocks_3_add_1_mdata_out_0;
assign fork2_8_edata_in_0 = stream_blocks_3_add_1_edata_out_0;

assign fork2_8_data_out_0_ready  = stream_blocks_4_linear1_data_in_0_ready;
assign stream_blocks_4_linear1_data_in_0_valid    = fork2_8_data_out_0_valid;
assign stream_blocks_4_linear1_mdata_in_0 = fork2_8_mdata_out_0;
assign stream_blocks_4_linear1_edata_in_0 = fork2_8_edata_out_0;

assign stream_blocks_4_linear1_data_out_0_ready  = stream_blocks_4_act_data_in_0_ready;
assign stream_blocks_4_act_data_in_0_valid    = stream_blocks_4_linear1_data_out_0_valid;
assign stream_blocks_4_act_mdata_in_0 = stream_blocks_4_linear1_mdata_out_0;
assign stream_blocks_4_act_edata_in_0 = stream_blocks_4_linear1_edata_out_0;

assign stream_blocks_4_act_data_out_0_ready  = stream_blocks_4_linear2_data_in_0_ready;
assign stream_blocks_4_linear2_data_in_0_valid    = stream_blocks_4_act_data_out_0_valid;
assign stream_blocks_4_linear2_mdata_in_0 = stream_blocks_4_act_mdata_out_0;
assign stream_blocks_4_linear2_edata_in_0 = stream_blocks_4_act_edata_out_0;

assign stream_blocks_4_linear2_data_out_0_ready  = stream_blocks_4_norm1_data_in_0_ready;
assign stream_blocks_4_norm1_data_in_0_valid    = stream_blocks_4_linear2_data_out_0_valid;
assign stream_blocks_4_norm1_mdata_in_0 = stream_blocks_4_linear2_mdata_out_0;
assign stream_blocks_4_norm1_edata_in_0 = stream_blocks_4_linear2_edata_out_0;

assign stream_blocks_4_norm1_data_out_0_ready  = stream_blocks_4_add_data_in_0_ready;
assign stream_blocks_4_add_data_in_0_valid    = stream_blocks_4_norm1_data_out_0_valid;
assign stream_blocks_4_add_mdata_in_0 = stream_blocks_4_norm1_mdata_out_0;
assign stream_blocks_4_add_edata_in_0 = stream_blocks_4_norm1_edata_out_0;

assign fork2_8_data_out_1_ready  = stream_blocks_4_add_data_in_1_ready;
assign stream_blocks_4_add_data_in_1_valid    = fork2_8_data_out_1_valid;
assign stream_blocks_4_add_mdata_in_1 = fork2_8_mdata_out_1;
assign stream_blocks_4_add_edata_in_1 = fork2_8_edata_out_1;

assign stream_blocks_4_add_data_out_0_ready  = fork2_9_data_in_0_ready;
assign fork2_9_data_in_0_valid    = stream_blocks_4_add_data_out_0_valid;
assign fork2_9_mdata_in_0 = stream_blocks_4_add_mdata_out_0;
assign fork2_9_edata_in_0 = stream_blocks_4_add_edata_out_0;

assign fork2_9_data_out_0_ready  = stream_blocks_4_attention_data_in_0_ready;
assign stream_blocks_4_attention_data_in_0_valid    = fork2_9_data_out_0_valid;
assign stream_blocks_4_attention_mdata_in_0 = fork2_9_mdata_out_0;
assign stream_blocks_4_attention_edata_in_0 = fork2_9_edata_out_0;

assign stream_blocks_4_attention_data_out_0_ready  = stream_blocks_4_norm2_data_in_0_ready;
assign stream_blocks_4_norm2_data_in_0_valid    = stream_blocks_4_attention_data_out_0_valid;
assign stream_blocks_4_norm2_mdata_in_0 = stream_blocks_4_attention_mdata_out_0;
assign stream_blocks_4_norm2_edata_in_0 = stream_blocks_4_attention_edata_out_0;

assign stream_blocks_4_norm2_data_out_0_ready  = stream_blocks_4_add_1_data_in_0_ready;
assign stream_blocks_4_add_1_data_in_0_valid    = stream_blocks_4_norm2_data_out_0_valid;
assign stream_blocks_4_add_1_mdata_in_0 = stream_blocks_4_norm2_mdata_out_0;
assign stream_blocks_4_add_1_edata_in_0 = stream_blocks_4_norm2_edata_out_0;

assign fork2_9_data_out_1_ready  = stream_blocks_4_add_1_data_in_1_ready;
assign stream_blocks_4_add_1_data_in_1_valid    = fork2_9_data_out_1_valid;
assign stream_blocks_4_add_1_mdata_in_1 = fork2_9_mdata_out_1;
assign stream_blocks_4_add_1_edata_in_1 = fork2_9_edata_out_1;

assign stream_blocks_4_add_1_data_out_0_ready  = fork2_10_data_in_0_ready;
assign fork2_10_data_in_0_valid    = stream_blocks_4_add_1_data_out_0_valid;
assign fork2_10_mdata_in_0 = stream_blocks_4_add_1_mdata_out_0;
assign fork2_10_edata_in_0 = stream_blocks_4_add_1_edata_out_0;

assign fork2_10_data_out_0_ready  = stream_blocks_5_linear1_data_in_0_ready;
assign stream_blocks_5_linear1_data_in_0_valid    = fork2_10_data_out_0_valid;
assign stream_blocks_5_linear1_mdata_in_0 = fork2_10_mdata_out_0;
assign stream_blocks_5_linear1_edata_in_0 = fork2_10_edata_out_0;

assign stream_blocks_5_linear1_data_out_0_ready  = stream_blocks_5_act_data_in_0_ready;
assign stream_blocks_5_act_data_in_0_valid    = stream_blocks_5_linear1_data_out_0_valid;
assign stream_blocks_5_act_mdata_in_0 = stream_blocks_5_linear1_mdata_out_0;
assign stream_blocks_5_act_edata_in_0 = stream_blocks_5_linear1_edata_out_0;

assign stream_blocks_5_act_data_out_0_ready  = stream_blocks_5_linear2_data_in_0_ready;
assign stream_blocks_5_linear2_data_in_0_valid    = stream_blocks_5_act_data_out_0_valid;
assign stream_blocks_5_linear2_mdata_in_0 = stream_blocks_5_act_mdata_out_0;
assign stream_blocks_5_linear2_edata_in_0 = stream_blocks_5_act_edata_out_0;

assign stream_blocks_5_linear2_data_out_0_ready  = stream_blocks_5_norm1_data_in_0_ready;
assign stream_blocks_5_norm1_data_in_0_valid    = stream_blocks_5_linear2_data_out_0_valid;
assign stream_blocks_5_norm1_mdata_in_0 = stream_blocks_5_linear2_mdata_out_0;
assign stream_blocks_5_norm1_edata_in_0 = stream_blocks_5_linear2_edata_out_0;

assign stream_blocks_5_norm1_data_out_0_ready  = stream_blocks_5_add_data_in_0_ready;
assign stream_blocks_5_add_data_in_0_valid    = stream_blocks_5_norm1_data_out_0_valid;
assign stream_blocks_5_add_mdata_in_0 = stream_blocks_5_norm1_mdata_out_0;
assign stream_blocks_5_add_edata_in_0 = stream_blocks_5_norm1_edata_out_0;

assign fork2_10_data_out_1_ready  = stream_blocks_5_add_data_in_1_ready;
assign stream_blocks_5_add_data_in_1_valid    = fork2_10_data_out_1_valid;
assign stream_blocks_5_add_mdata_in_1 = fork2_10_mdata_out_1;
assign stream_blocks_5_add_edata_in_1 = fork2_10_edata_out_1;

assign stream_blocks_5_add_data_out_0_ready  = fork2_11_data_in_0_ready;
assign fork2_11_data_in_0_valid    = stream_blocks_5_add_data_out_0_valid;
assign fork2_11_mdata_in_0 = stream_blocks_5_add_mdata_out_0;
assign fork2_11_edata_in_0 = stream_blocks_5_add_edata_out_0;

assign fork2_11_data_out_0_ready  = stream_blocks_5_attention_data_in_0_ready;
assign stream_blocks_5_attention_data_in_0_valid    = fork2_11_data_out_0_valid;
assign stream_blocks_5_attention_mdata_in_0 = fork2_11_mdata_out_0;
assign stream_blocks_5_attention_edata_in_0 = fork2_11_edata_out_0;

assign stream_blocks_5_attention_data_out_0_ready  = stream_blocks_5_norm2_data_in_0_ready;
assign stream_blocks_5_norm2_data_in_0_valid    = stream_blocks_5_attention_data_out_0_valid;
assign stream_blocks_5_norm2_mdata_in_0 = stream_blocks_5_attention_mdata_out_0;
assign stream_blocks_5_norm2_edata_in_0 = stream_blocks_5_attention_edata_out_0;

assign stream_blocks_5_norm2_data_out_0_ready  = stream_blocks_5_add_1_data_in_0_ready;
assign stream_blocks_5_add_1_data_in_0_valid    = stream_blocks_5_norm2_data_out_0_valid;
assign stream_blocks_5_add_1_mdata_in_0 = stream_blocks_5_norm2_mdata_out_0;
assign stream_blocks_5_add_1_edata_in_0 = stream_blocks_5_norm2_edata_out_0;

assign fork2_11_data_out_1_ready  = stream_blocks_5_add_1_data_in_1_ready;
assign stream_blocks_5_add_1_data_in_1_valid    = fork2_11_data_out_1_valid;
assign stream_blocks_5_add_1_mdata_in_1 = fork2_11_mdata_out_1;
assign stream_blocks_5_add_1_edata_in_1 = fork2_11_edata_out_1;

assign stream_blocks_5_add_1_data_out_0_ready  = fork2_12_data_in_0_ready;
assign fork2_12_data_in_0_valid    = stream_blocks_5_add_1_data_out_0_valid;
assign fork2_12_mdata_in_0 = stream_blocks_5_add_1_mdata_out_0;
assign fork2_12_edata_in_0 = stream_blocks_5_add_1_edata_out_0;

assign fork2_12_data_out_0_ready  = stream_blocks_6_linear1_data_in_0_ready;
assign stream_blocks_6_linear1_data_in_0_valid    = fork2_12_data_out_0_valid;
assign stream_blocks_6_linear1_mdata_in_0 = fork2_12_mdata_out_0;
assign stream_blocks_6_linear1_edata_in_0 = fork2_12_edata_out_0;

assign stream_blocks_6_linear1_data_out_0_ready  = stream_blocks_6_act_data_in_0_ready;
assign stream_blocks_6_act_data_in_0_valid    = stream_blocks_6_linear1_data_out_0_valid;
assign stream_blocks_6_act_mdata_in_0 = stream_blocks_6_linear1_mdata_out_0;
assign stream_blocks_6_act_edata_in_0 = stream_blocks_6_linear1_edata_out_0;

assign stream_blocks_6_act_data_out_0_ready  = stream_blocks_6_linear2_data_in_0_ready;
assign stream_blocks_6_linear2_data_in_0_valid    = stream_blocks_6_act_data_out_0_valid;
assign stream_blocks_6_linear2_mdata_in_0 = stream_blocks_6_act_mdata_out_0;
assign stream_blocks_6_linear2_edata_in_0 = stream_blocks_6_act_edata_out_0;

assign stream_blocks_6_linear2_data_out_0_ready  = stream_blocks_6_norm1_data_in_0_ready;
assign stream_blocks_6_norm1_data_in_0_valid    = stream_blocks_6_linear2_data_out_0_valid;
assign stream_blocks_6_norm1_mdata_in_0 = stream_blocks_6_linear2_mdata_out_0;
assign stream_blocks_6_norm1_edata_in_0 = stream_blocks_6_linear2_edata_out_0;

assign stream_blocks_6_norm1_data_out_0_ready  = stream_blocks_6_add_data_in_0_ready;
assign stream_blocks_6_add_data_in_0_valid    = stream_blocks_6_norm1_data_out_0_valid;
assign stream_blocks_6_add_mdata_in_0 = stream_blocks_6_norm1_mdata_out_0;
assign stream_blocks_6_add_edata_in_0 = stream_blocks_6_norm1_edata_out_0;

assign fork2_12_data_out_1_ready  = stream_blocks_6_add_data_in_1_ready;
assign stream_blocks_6_add_data_in_1_valid    = fork2_12_data_out_1_valid;
assign stream_blocks_6_add_mdata_in_1 = fork2_12_mdata_out_1;
assign stream_blocks_6_add_edata_in_1 = fork2_12_edata_out_1;

assign stream_blocks_6_add_data_out_0_ready  = fork2_13_data_in_0_ready;
assign fork2_13_data_in_0_valid    = stream_blocks_6_add_data_out_0_valid;
assign fork2_13_mdata_in_0 = stream_blocks_6_add_mdata_out_0;
assign fork2_13_edata_in_0 = stream_blocks_6_add_edata_out_0;

assign fork2_13_data_out_0_ready  = stream_blocks_6_attention_data_in_0_ready;
assign stream_blocks_6_attention_data_in_0_valid    = fork2_13_data_out_0_valid;
assign stream_blocks_6_attention_mdata_in_0 = fork2_13_mdata_out_0;
assign stream_blocks_6_attention_edata_in_0 = fork2_13_edata_out_0;

assign stream_blocks_6_attention_data_out_0_ready  = stream_blocks_6_norm2_data_in_0_ready;
assign stream_blocks_6_norm2_data_in_0_valid    = stream_blocks_6_attention_data_out_0_valid;
assign stream_blocks_6_norm2_mdata_in_0 = stream_blocks_6_attention_mdata_out_0;
assign stream_blocks_6_norm2_edata_in_0 = stream_blocks_6_attention_edata_out_0;

assign stream_blocks_6_norm2_data_out_0_ready  = stream_blocks_6_add_1_data_in_0_ready;
assign stream_blocks_6_add_1_data_in_0_valid    = stream_blocks_6_norm2_data_out_0_valid;
assign stream_blocks_6_add_1_mdata_in_0 = stream_blocks_6_norm2_mdata_out_0;
assign stream_blocks_6_add_1_edata_in_0 = stream_blocks_6_norm2_edata_out_0;

assign fork2_13_data_out_1_ready  = stream_blocks_6_add_1_data_in_1_ready;
assign stream_blocks_6_add_1_data_in_1_valid    = fork2_13_data_out_1_valid;
assign stream_blocks_6_add_1_mdata_in_1 = fork2_13_mdata_out_1;
assign stream_blocks_6_add_1_edata_in_1 = fork2_13_edata_out_1;

assign stream_blocks_6_add_1_data_out_0_ready  = fork2_14_data_in_0_ready;
assign fork2_14_data_in_0_valid    = stream_blocks_6_add_1_data_out_0_valid;
assign fork2_14_mdata_in_0 = stream_blocks_6_add_1_mdata_out_0;
assign fork2_14_edata_in_0 = stream_blocks_6_add_1_edata_out_0;

assign fork2_14_data_out_0_ready  = stream_blocks_7_linear1_data_in_0_ready;
assign stream_blocks_7_linear1_data_in_0_valid    = fork2_14_data_out_0_valid;
assign stream_blocks_7_linear1_mdata_in_0 = fork2_14_mdata_out_0;
assign stream_blocks_7_linear1_edata_in_0 = fork2_14_edata_out_0;

assign stream_blocks_7_linear1_data_out_0_ready  = stream_blocks_7_act_data_in_0_ready;
assign stream_blocks_7_act_data_in_0_valid    = stream_blocks_7_linear1_data_out_0_valid;
assign stream_blocks_7_act_mdata_in_0 = stream_blocks_7_linear1_mdata_out_0;
assign stream_blocks_7_act_edata_in_0 = stream_blocks_7_linear1_edata_out_0;

assign stream_blocks_7_act_data_out_0_ready  = stream_blocks_7_linear2_data_in_0_ready;
assign stream_blocks_7_linear2_data_in_0_valid    = stream_blocks_7_act_data_out_0_valid;
assign stream_blocks_7_linear2_mdata_in_0 = stream_blocks_7_act_mdata_out_0;
assign stream_blocks_7_linear2_edata_in_0 = stream_blocks_7_act_edata_out_0;

assign stream_blocks_7_linear2_data_out_0_ready  = stream_blocks_7_norm1_data_in_0_ready;
assign stream_blocks_7_norm1_data_in_0_valid    = stream_blocks_7_linear2_data_out_0_valid;
assign stream_blocks_7_norm1_mdata_in_0 = stream_blocks_7_linear2_mdata_out_0;
assign stream_blocks_7_norm1_edata_in_0 = stream_blocks_7_linear2_edata_out_0;

assign stream_blocks_7_norm1_data_out_0_ready  = stream_blocks_7_add_data_in_0_ready;
assign stream_blocks_7_add_data_in_0_valid    = stream_blocks_7_norm1_data_out_0_valid;
assign stream_blocks_7_add_mdata_in_0 = stream_blocks_7_norm1_mdata_out_0;
assign stream_blocks_7_add_edata_in_0 = stream_blocks_7_norm1_edata_out_0;

assign fork2_14_data_out_1_ready  = stream_blocks_7_add_data_in_1_ready;
assign stream_blocks_7_add_data_in_1_valid    = fork2_14_data_out_1_valid;
assign stream_blocks_7_add_mdata_in_1 = fork2_14_mdata_out_1;
assign stream_blocks_7_add_edata_in_1 = fork2_14_edata_out_1;

assign stream_blocks_7_add_data_out_0_ready  = fork2_15_data_in_0_ready;
assign fork2_15_data_in_0_valid    = stream_blocks_7_add_data_out_0_valid;
assign fork2_15_mdata_in_0 = stream_blocks_7_add_mdata_out_0;
assign fork2_15_edata_in_0 = stream_blocks_7_add_edata_out_0;

assign fork2_15_data_out_0_ready  = stream_blocks_7_attention_data_in_0_ready;
assign stream_blocks_7_attention_data_in_0_valid    = fork2_15_data_out_0_valid;
assign stream_blocks_7_attention_mdata_in_0 = fork2_15_mdata_out_0;
assign stream_blocks_7_attention_edata_in_0 = fork2_15_edata_out_0;

assign stream_blocks_7_attention_data_out_0_ready  = stream_blocks_7_norm2_data_in_0_ready;
assign stream_blocks_7_norm2_data_in_0_valid    = stream_blocks_7_attention_data_out_0_valid;
assign stream_blocks_7_norm2_mdata_in_0 = stream_blocks_7_attention_mdata_out_0;
assign stream_blocks_7_norm2_edata_in_0 = stream_blocks_7_attention_edata_out_0;

assign stream_blocks_7_norm2_data_out_0_ready  = stream_blocks_7_add_1_data_in_0_ready;
assign stream_blocks_7_add_1_data_in_0_valid    = stream_blocks_7_norm2_data_out_0_valid;
assign stream_blocks_7_add_1_mdata_in_0 = stream_blocks_7_norm2_mdata_out_0;
assign stream_blocks_7_add_1_edata_in_0 = stream_blocks_7_norm2_edata_out_0;

assign fork2_15_data_out_1_ready  = stream_blocks_7_add_1_data_in_1_ready;
assign stream_blocks_7_add_1_data_in_1_valid    = fork2_15_data_out_1_valid;
assign stream_blocks_7_add_1_mdata_in_1 = fork2_15_mdata_out_1;
assign stream_blocks_7_add_1_edata_in_1 = fork2_15_edata_out_1;

assign stream_blocks_7_add_1_data_out_0_ready  = fork2_16_data_in_0_ready;
assign fork2_16_data_in_0_valid    = stream_blocks_7_add_1_data_out_0_valid;
assign fork2_16_mdata_in_0 = stream_blocks_7_add_1_mdata_out_0;
assign fork2_16_edata_in_0 = stream_blocks_7_add_1_edata_out_0;

assign fork2_16_data_out_0_ready  = stream_blocks_8_linear1_data_in_0_ready;
assign stream_blocks_8_linear1_data_in_0_valid    = fork2_16_data_out_0_valid;
assign stream_blocks_8_linear1_mdata_in_0 = fork2_16_mdata_out_0;
assign stream_blocks_8_linear1_edata_in_0 = fork2_16_edata_out_0;

assign stream_blocks_8_linear1_data_out_0_ready  = stream_blocks_8_act_data_in_0_ready;
assign stream_blocks_8_act_data_in_0_valid    = stream_blocks_8_linear1_data_out_0_valid;
assign stream_blocks_8_act_mdata_in_0 = stream_blocks_8_linear1_mdata_out_0;
assign stream_blocks_8_act_edata_in_0 = stream_blocks_8_linear1_edata_out_0;

assign stream_blocks_8_act_data_out_0_ready  = stream_blocks_8_linear2_data_in_0_ready;
assign stream_blocks_8_linear2_data_in_0_valid    = stream_blocks_8_act_data_out_0_valid;
assign stream_blocks_8_linear2_mdata_in_0 = stream_blocks_8_act_mdata_out_0;
assign stream_blocks_8_linear2_edata_in_0 = stream_blocks_8_act_edata_out_0;

assign stream_blocks_8_linear2_data_out_0_ready  = stream_blocks_8_norm1_data_in_0_ready;
assign stream_blocks_8_norm1_data_in_0_valid    = stream_blocks_8_linear2_data_out_0_valid;
assign stream_blocks_8_norm1_mdata_in_0 = stream_blocks_8_linear2_mdata_out_0;
assign stream_blocks_8_norm1_edata_in_0 = stream_blocks_8_linear2_edata_out_0;

assign stream_blocks_8_norm1_data_out_0_ready  = stream_blocks_8_add_data_in_0_ready;
assign stream_blocks_8_add_data_in_0_valid    = stream_blocks_8_norm1_data_out_0_valid;
assign stream_blocks_8_add_mdata_in_0 = stream_blocks_8_norm1_mdata_out_0;
assign stream_blocks_8_add_edata_in_0 = stream_blocks_8_norm1_edata_out_0;

assign fork2_16_data_out_1_ready  = stream_blocks_8_add_data_in_1_ready;
assign stream_blocks_8_add_data_in_1_valid    = fork2_16_data_out_1_valid;
assign stream_blocks_8_add_mdata_in_1 = fork2_16_mdata_out_1;
assign stream_blocks_8_add_edata_in_1 = fork2_16_edata_out_1;

assign stream_blocks_8_add_data_out_0_ready  = fork2_17_data_in_0_ready;
assign fork2_17_data_in_0_valid    = stream_blocks_8_add_data_out_0_valid;
assign fork2_17_mdata_in_0 = stream_blocks_8_add_mdata_out_0;
assign fork2_17_edata_in_0 = stream_blocks_8_add_edata_out_0;

assign fork2_17_data_out_0_ready  = stream_blocks_8_attention_data_in_0_ready;
assign stream_blocks_8_attention_data_in_0_valid    = fork2_17_data_out_0_valid;
assign stream_blocks_8_attention_mdata_in_0 = fork2_17_mdata_out_0;
assign stream_blocks_8_attention_edata_in_0 = fork2_17_edata_out_0;

assign stream_blocks_8_attention_data_out_0_ready  = stream_blocks_8_norm2_data_in_0_ready;
assign stream_blocks_8_norm2_data_in_0_valid    = stream_blocks_8_attention_data_out_0_valid;
assign stream_blocks_8_norm2_mdata_in_0 = stream_blocks_8_attention_mdata_out_0;
assign stream_blocks_8_norm2_edata_in_0 = stream_blocks_8_attention_edata_out_0;

assign stream_blocks_8_norm2_data_out_0_ready  = stream_blocks_8_add_1_data_in_0_ready;
assign stream_blocks_8_add_1_data_in_0_valid    = stream_blocks_8_norm2_data_out_0_valid;
assign stream_blocks_8_add_1_mdata_in_0 = stream_blocks_8_norm2_mdata_out_0;
assign stream_blocks_8_add_1_edata_in_0 = stream_blocks_8_norm2_edata_out_0;

assign fork2_17_data_out_1_ready  = stream_blocks_8_add_1_data_in_1_ready;
assign stream_blocks_8_add_1_data_in_1_valid    = fork2_17_data_out_1_valid;
assign stream_blocks_8_add_1_mdata_in_1 = fork2_17_mdata_out_1;
assign stream_blocks_8_add_1_edata_in_1 = fork2_17_edata_out_1;

assign stream_blocks_8_add_1_data_out_0_ready  = fork2_18_data_in_0_ready;
assign fork2_18_data_in_0_valid    = stream_blocks_8_add_1_data_out_0_valid;
assign fork2_18_mdata_in_0 = stream_blocks_8_add_1_mdata_out_0;
assign fork2_18_edata_in_0 = stream_blocks_8_add_1_edata_out_0;

assign fork2_18_data_out_0_ready  = stream_blocks_9_linear1_data_in_0_ready;
assign stream_blocks_9_linear1_data_in_0_valid    = fork2_18_data_out_0_valid;
assign stream_blocks_9_linear1_mdata_in_0 = fork2_18_mdata_out_0;
assign stream_blocks_9_linear1_edata_in_0 = fork2_18_edata_out_0;

assign stream_blocks_9_linear1_data_out_0_ready  = stream_blocks_9_act_data_in_0_ready;
assign stream_blocks_9_act_data_in_0_valid    = stream_blocks_9_linear1_data_out_0_valid;
assign stream_blocks_9_act_mdata_in_0 = stream_blocks_9_linear1_mdata_out_0;
assign stream_blocks_9_act_edata_in_0 = stream_blocks_9_linear1_edata_out_0;

assign stream_blocks_9_act_data_out_0_ready  = stream_blocks_9_linear2_data_in_0_ready;
assign stream_blocks_9_linear2_data_in_0_valid    = stream_blocks_9_act_data_out_0_valid;
assign stream_blocks_9_linear2_mdata_in_0 = stream_blocks_9_act_mdata_out_0;
assign stream_blocks_9_linear2_edata_in_0 = stream_blocks_9_act_edata_out_0;

assign stream_blocks_9_linear2_data_out_0_ready  = stream_blocks_9_norm1_data_in_0_ready;
assign stream_blocks_9_norm1_data_in_0_valid    = stream_blocks_9_linear2_data_out_0_valid;
assign stream_blocks_9_norm1_mdata_in_0 = stream_blocks_9_linear2_mdata_out_0;
assign stream_blocks_9_norm1_edata_in_0 = stream_blocks_9_linear2_edata_out_0;

assign stream_blocks_9_norm1_data_out_0_ready  = stream_blocks_9_add_data_in_0_ready;
assign stream_blocks_9_add_data_in_0_valid    = stream_blocks_9_norm1_data_out_0_valid;
assign stream_blocks_9_add_mdata_in_0 = stream_blocks_9_norm1_mdata_out_0;
assign stream_blocks_9_add_edata_in_0 = stream_blocks_9_norm1_edata_out_0;

assign fork2_18_data_out_1_ready  = stream_blocks_9_add_data_in_1_ready;
assign stream_blocks_9_add_data_in_1_valid    = fork2_18_data_out_1_valid;
assign stream_blocks_9_add_mdata_in_1 = fork2_18_mdata_out_1;
assign stream_blocks_9_add_edata_in_1 = fork2_18_edata_out_1;

assign stream_blocks_9_add_data_out_0_ready  = fork2_19_data_in_0_ready;
assign fork2_19_data_in_0_valid    = stream_blocks_9_add_data_out_0_valid;
assign fork2_19_mdata_in_0 = stream_blocks_9_add_mdata_out_0;
assign fork2_19_edata_in_0 = stream_blocks_9_add_edata_out_0;

assign fork2_19_data_out_0_ready  = stream_blocks_9_attention_data_in_0_ready;
assign stream_blocks_9_attention_data_in_0_valid    = fork2_19_data_out_0_valid;
assign stream_blocks_9_attention_mdata_in_0 = fork2_19_mdata_out_0;
assign stream_blocks_9_attention_edata_in_0 = fork2_19_edata_out_0;

assign stream_blocks_9_attention_data_out_0_ready  = stream_blocks_9_norm2_data_in_0_ready;
assign stream_blocks_9_norm2_data_in_0_valid    = stream_blocks_9_attention_data_out_0_valid;
assign stream_blocks_9_norm2_mdata_in_0 = stream_blocks_9_attention_mdata_out_0;
assign stream_blocks_9_norm2_edata_in_0 = stream_blocks_9_attention_edata_out_0;

assign stream_blocks_9_norm2_data_out_0_ready  = stream_blocks_9_add_1_data_in_0_ready;
assign stream_blocks_9_add_1_data_in_0_valid    = stream_blocks_9_norm2_data_out_0_valid;
assign stream_blocks_9_add_1_mdata_in_0 = stream_blocks_9_norm2_mdata_out_0;
assign stream_blocks_9_add_1_edata_in_0 = stream_blocks_9_norm2_edata_out_0;

assign fork2_19_data_out_1_ready  = stream_blocks_9_add_1_data_in_1_ready;
assign stream_blocks_9_add_1_data_in_1_valid    = fork2_19_data_out_1_valid;
assign stream_blocks_9_add_1_mdata_in_1 = fork2_19_mdata_out_1;
assign stream_blocks_9_add_1_edata_in_1 = fork2_19_edata_out_1;

assign stream_blocks_9_add_1_data_out_0_ready  = fork2_20_data_in_0_ready;
assign fork2_20_data_in_0_valid    = stream_blocks_9_add_1_data_out_0_valid;
assign fork2_20_mdata_in_0 = stream_blocks_9_add_1_mdata_out_0;
assign fork2_20_edata_in_0 = stream_blocks_9_add_1_edata_out_0;

assign fork2_20_data_out_0_ready  = stream_blocks_10_linear1_data_in_0_ready;
assign stream_blocks_10_linear1_data_in_0_valid    = fork2_20_data_out_0_valid;
assign stream_blocks_10_linear1_mdata_in_0 = fork2_20_mdata_out_0;
assign stream_blocks_10_linear1_edata_in_0 = fork2_20_edata_out_0;

assign stream_blocks_10_linear1_data_out_0_ready  = stream_blocks_10_act_data_in_0_ready;
assign stream_blocks_10_act_data_in_0_valid    = stream_blocks_10_linear1_data_out_0_valid;
assign stream_blocks_10_act_mdata_in_0 = stream_blocks_10_linear1_mdata_out_0;
assign stream_blocks_10_act_edata_in_0 = stream_blocks_10_linear1_edata_out_0;

assign stream_blocks_10_act_data_out_0_ready  = stream_blocks_10_linear2_data_in_0_ready;
assign stream_blocks_10_linear2_data_in_0_valid    = stream_blocks_10_act_data_out_0_valid;
assign stream_blocks_10_linear2_mdata_in_0 = stream_blocks_10_act_mdata_out_0;
assign stream_blocks_10_linear2_edata_in_0 = stream_blocks_10_act_edata_out_0;

assign stream_blocks_10_linear2_data_out_0_ready  = stream_blocks_10_norm1_data_in_0_ready;
assign stream_blocks_10_norm1_data_in_0_valid    = stream_blocks_10_linear2_data_out_0_valid;
assign stream_blocks_10_norm1_mdata_in_0 = stream_blocks_10_linear2_mdata_out_0;
assign stream_blocks_10_norm1_edata_in_0 = stream_blocks_10_linear2_edata_out_0;

assign stream_blocks_10_norm1_data_out_0_ready  = stream_blocks_10_add_data_in_0_ready;
assign stream_blocks_10_add_data_in_0_valid    = stream_blocks_10_norm1_data_out_0_valid;
assign stream_blocks_10_add_mdata_in_0 = stream_blocks_10_norm1_mdata_out_0;
assign stream_blocks_10_add_edata_in_0 = stream_blocks_10_norm1_edata_out_0;

assign fork2_20_data_out_1_ready  = stream_blocks_10_add_data_in_1_ready;
assign stream_blocks_10_add_data_in_1_valid    = fork2_20_data_out_1_valid;
assign stream_blocks_10_add_mdata_in_1 = fork2_20_mdata_out_1;
assign stream_blocks_10_add_edata_in_1 = fork2_20_edata_out_1;

assign stream_blocks_10_add_data_out_0_ready  = fork2_21_data_in_0_ready;
assign fork2_21_data_in_0_valid    = stream_blocks_10_add_data_out_0_valid;
assign fork2_21_mdata_in_0 = stream_blocks_10_add_mdata_out_0;
assign fork2_21_edata_in_0 = stream_blocks_10_add_edata_out_0;

assign fork2_21_data_out_0_ready  = stream_blocks_10_attention_data_in_0_ready;
assign stream_blocks_10_attention_data_in_0_valid    = fork2_21_data_out_0_valid;
assign stream_blocks_10_attention_mdata_in_0 = fork2_21_mdata_out_0;
assign stream_blocks_10_attention_edata_in_0 = fork2_21_edata_out_0;

assign stream_blocks_10_attention_data_out_0_ready  = stream_blocks_10_norm2_data_in_0_ready;
assign stream_blocks_10_norm2_data_in_0_valid    = stream_blocks_10_attention_data_out_0_valid;
assign stream_blocks_10_norm2_mdata_in_0 = stream_blocks_10_attention_mdata_out_0;
assign stream_blocks_10_norm2_edata_in_0 = stream_blocks_10_attention_edata_out_0;

assign stream_blocks_10_norm2_data_out_0_ready  = stream_blocks_10_add_1_data_in_0_ready;
assign stream_blocks_10_add_1_data_in_0_valid    = stream_blocks_10_norm2_data_out_0_valid;
assign stream_blocks_10_add_1_mdata_in_0 = stream_blocks_10_norm2_mdata_out_0;
assign stream_blocks_10_add_1_edata_in_0 = stream_blocks_10_norm2_edata_out_0;

assign fork2_21_data_out_1_ready  = stream_blocks_10_add_1_data_in_1_ready;
assign stream_blocks_10_add_1_data_in_1_valid    = fork2_21_data_out_1_valid;
assign stream_blocks_10_add_1_mdata_in_1 = fork2_21_mdata_out_1;
assign stream_blocks_10_add_1_edata_in_1 = fork2_21_edata_out_1;

assign stream_blocks_10_add_1_data_out_0_ready  = fork2_22_data_in_0_ready;
assign fork2_22_data_in_0_valid    = stream_blocks_10_add_1_data_out_0_valid;
assign fork2_22_mdata_in_0 = stream_blocks_10_add_1_mdata_out_0;
assign fork2_22_edata_in_0 = stream_blocks_10_add_1_edata_out_0;

assign fork2_22_data_out_0_ready  = stream_blocks_11_linear1_data_in_0_ready;
assign stream_blocks_11_linear1_data_in_0_valid    = fork2_22_data_out_0_valid;
assign stream_blocks_11_linear1_mdata_in_0 = fork2_22_mdata_out_0;
assign stream_blocks_11_linear1_edata_in_0 = fork2_22_edata_out_0;

assign stream_blocks_11_linear1_data_out_0_ready  = stream_blocks_11_act_data_in_0_ready;
assign stream_blocks_11_act_data_in_0_valid    = stream_blocks_11_linear1_data_out_0_valid;
assign stream_blocks_11_act_mdata_in_0 = stream_blocks_11_linear1_mdata_out_0;
assign stream_blocks_11_act_edata_in_0 = stream_blocks_11_linear1_edata_out_0;

assign stream_blocks_11_act_data_out_0_ready  = stream_blocks_11_linear2_data_in_0_ready;
assign stream_blocks_11_linear2_data_in_0_valid    = stream_blocks_11_act_data_out_0_valid;
assign stream_blocks_11_linear2_mdata_in_0 = stream_blocks_11_act_mdata_out_0;
assign stream_blocks_11_linear2_edata_in_0 = stream_blocks_11_act_edata_out_0;

assign stream_blocks_11_linear2_data_out_0_ready  = stream_blocks_11_norm1_data_in_0_ready;
assign stream_blocks_11_norm1_data_in_0_valid    = stream_blocks_11_linear2_data_out_0_valid;
assign stream_blocks_11_norm1_mdata_in_0 = stream_blocks_11_linear2_mdata_out_0;
assign stream_blocks_11_norm1_edata_in_0 = stream_blocks_11_linear2_edata_out_0;

assign stream_blocks_11_norm1_data_out_0_ready  = stream_blocks_11_add_data_in_0_ready;
assign stream_blocks_11_add_data_in_0_valid    = stream_blocks_11_norm1_data_out_0_valid;
assign stream_blocks_11_add_mdata_in_0 = stream_blocks_11_norm1_mdata_out_0;
assign stream_blocks_11_add_edata_in_0 = stream_blocks_11_norm1_edata_out_0;

assign fork2_22_data_out_1_ready  = stream_blocks_11_add_data_in_1_ready;
assign stream_blocks_11_add_data_in_1_valid    = fork2_22_data_out_1_valid;
assign stream_blocks_11_add_mdata_in_1 = fork2_22_mdata_out_1;
assign stream_blocks_11_add_edata_in_1 = fork2_22_edata_out_1;

assign stream_blocks_11_add_data_out_0_ready  = fork2_23_data_in_0_ready;
assign fork2_23_data_in_0_valid    = stream_blocks_11_add_data_out_0_valid;
assign fork2_23_mdata_in_0 = stream_blocks_11_add_mdata_out_0;
assign fork2_23_edata_in_0 = stream_blocks_11_add_edata_out_0;

assign fork2_23_data_out_0_ready  = stream_blocks_11_attention_data_in_0_ready;
assign stream_blocks_11_attention_data_in_0_valid    = fork2_23_data_out_0_valid;
assign stream_blocks_11_attention_mdata_in_0 = fork2_23_mdata_out_0;
assign stream_blocks_11_attention_edata_in_0 = fork2_23_edata_out_0;

assign stream_blocks_11_attention_data_out_0_ready  = stream_blocks_11_norm2_data_in_0_ready;
assign stream_blocks_11_norm2_data_in_0_valid    = stream_blocks_11_attention_data_out_0_valid;
assign stream_blocks_11_norm2_mdata_in_0 = stream_blocks_11_attention_mdata_out_0;
assign stream_blocks_11_norm2_edata_in_0 = stream_blocks_11_attention_edata_out_0;

assign stream_blocks_11_norm2_data_out_0_ready  = stream_blocks_11_add_1_data_in_0_ready;
assign stream_blocks_11_add_1_data_in_0_valid    = stream_blocks_11_norm2_data_out_0_valid;
assign stream_blocks_11_add_1_mdata_in_0 = stream_blocks_11_norm2_mdata_out_0;
assign stream_blocks_11_add_1_edata_in_0 = stream_blocks_11_norm2_edata_out_0;

assign fork2_23_data_out_1_ready  = stream_blocks_11_add_1_data_in_1_ready;
assign stream_blocks_11_add_1_data_in_1_valid    = fork2_23_data_out_1_valid;
assign stream_blocks_11_add_1_mdata_in_1 = fork2_23_mdata_out_1;
assign stream_blocks_11_add_1_edata_in_1 = fork2_23_edata_out_1;

endmodule
    
    
`timescale 1ns / 1ps
module stream_blocks_0_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_linear1_eweight;
logic folded_blocks_0_stream_blocks_0_linear1_weight_valid, folded_blocks_0_stream_blocks_0_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_0_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_0_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear1_mweight: folded_blocks_0_stream_blocks_0_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear1_eweight: folded_blocks_0_stream_blocks_0_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear1_weight_valid: folded_blocks_0_stream_blocks_0_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_linear1_ebias;
logic folded_blocks_0_stream_blocks_0_linear1_bias_valid, folded_blocks_0_stream_blocks_0_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_0_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_0_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear1_mbias: folded_blocks_0_stream_blocks_0_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear1_ebias: folded_blocks_0_stream_blocks_0_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear1_bias_valid: folded_blocks_0_stream_blocks_0_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_linear2_eweight;
logic folded_blocks_0_stream_blocks_0_linear2_weight_valid, folded_blocks_0_stream_blocks_0_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_0_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_0_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear2_mweight: folded_blocks_0_stream_blocks_0_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear2_eweight: folded_blocks_0_stream_blocks_0_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear2_weight_valid: folded_blocks_0_stream_blocks_0_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_linear2_ebias;
logic folded_blocks_0_stream_blocks_0_linear2_bias_valid, folded_blocks_0_stream_blocks_0_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_0_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_0_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear2_mbias: folded_blocks_0_stream_blocks_0_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear2_ebias: folded_blocks_0_stream_blocks_0_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_linear2_bias_valid: folded_blocks_0_stream_blocks_0_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_norm1_eweight;
logic folded_blocks_0_stream_blocks_0_norm1_weight_valid, folded_blocks_0_stream_blocks_0_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_0_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_0_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm1_mweight: folded_blocks_0_stream_blocks_0_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm1_eweight: folded_blocks_0_stream_blocks_0_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm1_weight_valid: folded_blocks_0_stream_blocks_0_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_norm1_ebias;
logic folded_blocks_0_stream_blocks_0_norm1_bias_valid, folded_blocks_0_stream_blocks_0_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_0_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_0_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm1_mbias: folded_blocks_0_stream_blocks_0_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm1_ebias: folded_blocks_0_stream_blocks_0_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm1_bias_valid: folded_blocks_0_stream_blocks_0_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_attention_equery_weight;
logic folded_blocks_0_stream_blocks_0_attention_query_weight_valid, folded_blocks_0_stream_blocks_0_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_0_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_0_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_mquery_weight: folded_blocks_0_stream_blocks_0_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_equery_weight: folded_blocks_0_stream_blocks_0_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_query_weight_valid: folded_blocks_0_stream_blocks_0_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_attention_equery_bias;
logic folded_blocks_0_stream_blocks_0_attention_query_bias_valid, folded_blocks_0_stream_blocks_0_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_0_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_0_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_mquery_bias: folded_blocks_0_stream_blocks_0_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_equery_bias: folded_blocks_0_stream_blocks_0_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_query_bias_valid: folded_blocks_0_stream_blocks_0_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_0_attention_key_weight_valid, folded_blocks_0_stream_blocks_0_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_0_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_0_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_mkey_weight: folded_blocks_0_stream_blocks_0_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_ekey_weight: folded_blocks_0_stream_blocks_0_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_key_weight_valid: folded_blocks_0_stream_blocks_0_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_0_attention_key_bias_valid, folded_blocks_0_stream_blocks_0_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_0_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_0_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_mkey_bias: folded_blocks_0_stream_blocks_0_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_ekey_bias: folded_blocks_0_stream_blocks_0_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_key_bias_valid: folded_blocks_0_stream_blocks_0_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_0_attention_value_weight_valid, folded_blocks_0_stream_blocks_0_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_0_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_0_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_mvalue_weight: folded_blocks_0_stream_blocks_0_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_evalue_weight: folded_blocks_0_stream_blocks_0_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_value_weight_valid: folded_blocks_0_stream_blocks_0_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_0_attention_value_bias_valid, folded_blocks_0_stream_blocks_0_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_0_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_0_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_mvalue_bias: folded_blocks_0_stream_blocks_0_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_evalue_bias: folded_blocks_0_stream_blocks_0_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_value_bias_valid: folded_blocks_0_stream_blocks_0_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_0_attention_proj_weight_valid, folded_blocks_0_stream_blocks_0_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_0_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_0_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_mproj_weight: folded_blocks_0_stream_blocks_0_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_eproj_weight: folded_blocks_0_stream_blocks_0_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_proj_weight_valid: folded_blocks_0_stream_blocks_0_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_0_attention_proj_bias_valid, folded_blocks_0_stream_blocks_0_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_0_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_0_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_mproj_bias: folded_blocks_0_stream_blocks_0_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_eproj_bias: folded_blocks_0_stream_blocks_0_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_attention_proj_bias_valid: folded_blocks_0_stream_blocks_0_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_norm2_eweight;
logic folded_blocks_0_stream_blocks_0_norm2_weight_valid, folded_blocks_0_stream_blocks_0_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_0_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_0_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm2_mweight: folded_blocks_0_stream_blocks_0_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm2_eweight: folded_blocks_0_stream_blocks_0_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm2_weight_valid: folded_blocks_0_stream_blocks_0_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_0_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_0_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_0_norm2_ebias;
logic folded_blocks_0_stream_blocks_0_norm2_bias_valid, folded_blocks_0_stream_blocks_0_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_0_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_0_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_0_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_0_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_0_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_0_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_0_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm2_mbias: folded_blocks_0_stream_blocks_0_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm2_ebias: folded_blocks_0_stream_blocks_0_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_0_norm2_bias_valid: folded_blocks_0_stream_blocks_0_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_linear1_eweight;
logic folded_blocks_0_stream_blocks_1_linear1_weight_valid, folded_blocks_0_stream_blocks_1_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_1_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_1_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear1_mweight: folded_blocks_0_stream_blocks_1_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear1_eweight: folded_blocks_0_stream_blocks_1_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear1_weight_valid: folded_blocks_0_stream_blocks_1_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_linear1_ebias;
logic folded_blocks_0_stream_blocks_1_linear1_bias_valid, folded_blocks_0_stream_blocks_1_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_1_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_1_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear1_mbias: folded_blocks_0_stream_blocks_1_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear1_ebias: folded_blocks_0_stream_blocks_1_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear1_bias_valid: folded_blocks_0_stream_blocks_1_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_linear2_eweight;
logic folded_blocks_0_stream_blocks_1_linear2_weight_valid, folded_blocks_0_stream_blocks_1_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_1_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_1_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear2_mweight: folded_blocks_0_stream_blocks_1_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear2_eweight: folded_blocks_0_stream_blocks_1_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear2_weight_valid: folded_blocks_0_stream_blocks_1_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_linear2_ebias;
logic folded_blocks_0_stream_blocks_1_linear2_bias_valid, folded_blocks_0_stream_blocks_1_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_1_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_1_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear2_mbias: folded_blocks_0_stream_blocks_1_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear2_ebias: folded_blocks_0_stream_blocks_1_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_linear2_bias_valid: folded_blocks_0_stream_blocks_1_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_norm1_eweight;
logic folded_blocks_0_stream_blocks_1_norm1_weight_valid, folded_blocks_0_stream_blocks_1_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_1_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_1_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm1_mweight: folded_blocks_0_stream_blocks_1_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm1_eweight: folded_blocks_0_stream_blocks_1_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm1_weight_valid: folded_blocks_0_stream_blocks_1_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_norm1_ebias;
logic folded_blocks_0_stream_blocks_1_norm1_bias_valid, folded_blocks_0_stream_blocks_1_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_1_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_1_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm1_mbias: folded_blocks_0_stream_blocks_1_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm1_ebias: folded_blocks_0_stream_blocks_1_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm1_bias_valid: folded_blocks_0_stream_blocks_1_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_attention_equery_weight;
logic folded_blocks_0_stream_blocks_1_attention_query_weight_valid, folded_blocks_0_stream_blocks_1_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_1_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_1_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_mquery_weight: folded_blocks_0_stream_blocks_1_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_equery_weight: folded_blocks_0_stream_blocks_1_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_query_weight_valid: folded_blocks_0_stream_blocks_1_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_attention_equery_bias;
logic folded_blocks_0_stream_blocks_1_attention_query_bias_valid, folded_blocks_0_stream_blocks_1_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_1_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_1_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_mquery_bias: folded_blocks_0_stream_blocks_1_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_equery_bias: folded_blocks_0_stream_blocks_1_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_query_bias_valid: folded_blocks_0_stream_blocks_1_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_1_attention_key_weight_valid, folded_blocks_0_stream_blocks_1_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_1_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_1_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_mkey_weight: folded_blocks_0_stream_blocks_1_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_ekey_weight: folded_blocks_0_stream_blocks_1_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_key_weight_valid: folded_blocks_0_stream_blocks_1_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_1_attention_key_bias_valid, folded_blocks_0_stream_blocks_1_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_1_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_1_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_mkey_bias: folded_blocks_0_stream_blocks_1_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_ekey_bias: folded_blocks_0_stream_blocks_1_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_key_bias_valid: folded_blocks_0_stream_blocks_1_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_1_attention_value_weight_valid, folded_blocks_0_stream_blocks_1_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_1_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_1_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_mvalue_weight: folded_blocks_0_stream_blocks_1_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_evalue_weight: folded_blocks_0_stream_blocks_1_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_value_weight_valid: folded_blocks_0_stream_blocks_1_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_1_attention_value_bias_valid, folded_blocks_0_stream_blocks_1_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_1_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_1_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_mvalue_bias: folded_blocks_0_stream_blocks_1_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_evalue_bias: folded_blocks_0_stream_blocks_1_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_value_bias_valid: folded_blocks_0_stream_blocks_1_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_1_attention_proj_weight_valid, folded_blocks_0_stream_blocks_1_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_1_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_1_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_mproj_weight: folded_blocks_0_stream_blocks_1_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_eproj_weight: folded_blocks_0_stream_blocks_1_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_proj_weight_valid: folded_blocks_0_stream_blocks_1_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_1_attention_proj_bias_valid, folded_blocks_0_stream_blocks_1_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_1_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_1_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_mproj_bias: folded_blocks_0_stream_blocks_1_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_eproj_bias: folded_blocks_0_stream_blocks_1_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_attention_proj_bias_valid: folded_blocks_0_stream_blocks_1_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_norm2_eweight;
logic folded_blocks_0_stream_blocks_1_norm2_weight_valid, folded_blocks_0_stream_blocks_1_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_1_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_1_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm2_mweight: folded_blocks_0_stream_blocks_1_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm2_eweight: folded_blocks_0_stream_blocks_1_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm2_weight_valid: folded_blocks_0_stream_blocks_1_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_1_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_1_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_1_norm2_ebias;
logic folded_blocks_0_stream_blocks_1_norm2_bias_valid, folded_blocks_0_stream_blocks_1_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_1_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_1_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_1_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_1_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_1_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_1_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_1_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm2_mbias: folded_blocks_0_stream_blocks_1_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm2_ebias: folded_blocks_0_stream_blocks_1_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_1_norm2_bias_valid: folded_blocks_0_stream_blocks_1_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_linear1_eweight;
logic folded_blocks_0_stream_blocks_2_linear1_weight_valid, folded_blocks_0_stream_blocks_2_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_2_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_2_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear1_mweight: folded_blocks_0_stream_blocks_2_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear1_eweight: folded_blocks_0_stream_blocks_2_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear1_weight_valid: folded_blocks_0_stream_blocks_2_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_linear1_ebias;
logic folded_blocks_0_stream_blocks_2_linear1_bias_valid, folded_blocks_0_stream_blocks_2_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_2_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_2_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear1_mbias: folded_blocks_0_stream_blocks_2_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear1_ebias: folded_blocks_0_stream_blocks_2_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear1_bias_valid: folded_blocks_0_stream_blocks_2_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_linear2_eweight;
logic folded_blocks_0_stream_blocks_2_linear2_weight_valid, folded_blocks_0_stream_blocks_2_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_2_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_2_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear2_mweight: folded_blocks_0_stream_blocks_2_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear2_eweight: folded_blocks_0_stream_blocks_2_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear2_weight_valid: folded_blocks_0_stream_blocks_2_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_linear2_ebias;
logic folded_blocks_0_stream_blocks_2_linear2_bias_valid, folded_blocks_0_stream_blocks_2_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_2_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_2_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear2_mbias: folded_blocks_0_stream_blocks_2_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear2_ebias: folded_blocks_0_stream_blocks_2_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_linear2_bias_valid: folded_blocks_0_stream_blocks_2_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_norm1_eweight;
logic folded_blocks_0_stream_blocks_2_norm1_weight_valid, folded_blocks_0_stream_blocks_2_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_2_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_2_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm1_mweight: folded_blocks_0_stream_blocks_2_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm1_eweight: folded_blocks_0_stream_blocks_2_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm1_weight_valid: folded_blocks_0_stream_blocks_2_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_norm1_ebias;
logic folded_blocks_0_stream_blocks_2_norm1_bias_valid, folded_blocks_0_stream_blocks_2_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_2_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_2_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm1_mbias: folded_blocks_0_stream_blocks_2_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm1_ebias: folded_blocks_0_stream_blocks_2_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm1_bias_valid: folded_blocks_0_stream_blocks_2_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_attention_equery_weight;
logic folded_blocks_0_stream_blocks_2_attention_query_weight_valid, folded_blocks_0_stream_blocks_2_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_2_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_2_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_mquery_weight: folded_blocks_0_stream_blocks_2_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_equery_weight: folded_blocks_0_stream_blocks_2_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_query_weight_valid: folded_blocks_0_stream_blocks_2_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_attention_equery_bias;
logic folded_blocks_0_stream_blocks_2_attention_query_bias_valid, folded_blocks_0_stream_blocks_2_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_2_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_2_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_mquery_bias: folded_blocks_0_stream_blocks_2_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_equery_bias: folded_blocks_0_stream_blocks_2_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_query_bias_valid: folded_blocks_0_stream_blocks_2_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_2_attention_key_weight_valid, folded_blocks_0_stream_blocks_2_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_2_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_2_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_mkey_weight: folded_blocks_0_stream_blocks_2_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_ekey_weight: folded_blocks_0_stream_blocks_2_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_key_weight_valid: folded_blocks_0_stream_blocks_2_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_2_attention_key_bias_valid, folded_blocks_0_stream_blocks_2_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_2_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_2_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_mkey_bias: folded_blocks_0_stream_blocks_2_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_ekey_bias: folded_blocks_0_stream_blocks_2_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_key_bias_valid: folded_blocks_0_stream_blocks_2_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_2_attention_value_weight_valid, folded_blocks_0_stream_blocks_2_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_2_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_2_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_mvalue_weight: folded_blocks_0_stream_blocks_2_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_evalue_weight: folded_blocks_0_stream_blocks_2_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_value_weight_valid: folded_blocks_0_stream_blocks_2_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_2_attention_value_bias_valid, folded_blocks_0_stream_blocks_2_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_2_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_2_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_mvalue_bias: folded_blocks_0_stream_blocks_2_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_evalue_bias: folded_blocks_0_stream_blocks_2_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_value_bias_valid: folded_blocks_0_stream_blocks_2_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_2_attention_proj_weight_valid, folded_blocks_0_stream_blocks_2_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_2_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_2_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_mproj_weight: folded_blocks_0_stream_blocks_2_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_eproj_weight: folded_blocks_0_stream_blocks_2_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_proj_weight_valid: folded_blocks_0_stream_blocks_2_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_2_attention_proj_bias_valid, folded_blocks_0_stream_blocks_2_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_2_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_2_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_mproj_bias: folded_blocks_0_stream_blocks_2_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_eproj_bias: folded_blocks_0_stream_blocks_2_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_attention_proj_bias_valid: folded_blocks_0_stream_blocks_2_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_norm2_eweight;
logic folded_blocks_0_stream_blocks_2_norm2_weight_valid, folded_blocks_0_stream_blocks_2_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_2_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_2_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm2_mweight: folded_blocks_0_stream_blocks_2_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm2_eweight: folded_blocks_0_stream_blocks_2_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm2_weight_valid: folded_blocks_0_stream_blocks_2_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_2_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_2_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_2_norm2_ebias;
logic folded_blocks_0_stream_blocks_2_norm2_bias_valid, folded_blocks_0_stream_blocks_2_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_2_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_2_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_2_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_2_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_2_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_2_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_2_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm2_mbias: folded_blocks_0_stream_blocks_2_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm2_ebias: folded_blocks_0_stream_blocks_2_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_2_norm2_bias_valid: folded_blocks_0_stream_blocks_2_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_linear1_eweight;
logic folded_blocks_0_stream_blocks_3_linear1_weight_valid, folded_blocks_0_stream_blocks_3_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_3_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_3_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear1_mweight: folded_blocks_0_stream_blocks_3_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear1_eweight: folded_blocks_0_stream_blocks_3_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear1_weight_valid: folded_blocks_0_stream_blocks_3_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_linear1_ebias;
logic folded_blocks_0_stream_blocks_3_linear1_bias_valid, folded_blocks_0_stream_blocks_3_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_3_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_3_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear1_mbias: folded_blocks_0_stream_blocks_3_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear1_ebias: folded_blocks_0_stream_blocks_3_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear1_bias_valid: folded_blocks_0_stream_blocks_3_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_linear2_eweight;
logic folded_blocks_0_stream_blocks_3_linear2_weight_valid, folded_blocks_0_stream_blocks_3_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_3_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_3_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear2_mweight: folded_blocks_0_stream_blocks_3_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear2_eweight: folded_blocks_0_stream_blocks_3_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear2_weight_valid: folded_blocks_0_stream_blocks_3_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_linear2_ebias;
logic folded_blocks_0_stream_blocks_3_linear2_bias_valid, folded_blocks_0_stream_blocks_3_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_3_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_3_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear2_mbias: folded_blocks_0_stream_blocks_3_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear2_ebias: folded_blocks_0_stream_blocks_3_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_linear2_bias_valid: folded_blocks_0_stream_blocks_3_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_norm1_eweight;
logic folded_blocks_0_stream_blocks_3_norm1_weight_valid, folded_blocks_0_stream_blocks_3_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_3_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_3_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm1_mweight: folded_blocks_0_stream_blocks_3_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm1_eweight: folded_blocks_0_stream_blocks_3_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm1_weight_valid: folded_blocks_0_stream_blocks_3_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_norm1_ebias;
logic folded_blocks_0_stream_blocks_3_norm1_bias_valid, folded_blocks_0_stream_blocks_3_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_3_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_3_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm1_mbias: folded_blocks_0_stream_blocks_3_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm1_ebias: folded_blocks_0_stream_blocks_3_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm1_bias_valid: folded_blocks_0_stream_blocks_3_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_attention_equery_weight;
logic folded_blocks_0_stream_blocks_3_attention_query_weight_valid, folded_blocks_0_stream_blocks_3_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_3_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_3_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_mquery_weight: folded_blocks_0_stream_blocks_3_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_equery_weight: folded_blocks_0_stream_blocks_3_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_query_weight_valid: folded_blocks_0_stream_blocks_3_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_attention_equery_bias;
logic folded_blocks_0_stream_blocks_3_attention_query_bias_valid, folded_blocks_0_stream_blocks_3_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_3_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_3_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_mquery_bias: folded_blocks_0_stream_blocks_3_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_equery_bias: folded_blocks_0_stream_blocks_3_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_query_bias_valid: folded_blocks_0_stream_blocks_3_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_3_attention_key_weight_valid, folded_blocks_0_stream_blocks_3_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_3_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_3_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_mkey_weight: folded_blocks_0_stream_blocks_3_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_ekey_weight: folded_blocks_0_stream_blocks_3_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_key_weight_valid: folded_blocks_0_stream_blocks_3_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_3_attention_key_bias_valid, folded_blocks_0_stream_blocks_3_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_3_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_3_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_mkey_bias: folded_blocks_0_stream_blocks_3_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_ekey_bias: folded_blocks_0_stream_blocks_3_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_key_bias_valid: folded_blocks_0_stream_blocks_3_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_3_attention_value_weight_valid, folded_blocks_0_stream_blocks_3_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_3_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_3_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_mvalue_weight: folded_blocks_0_stream_blocks_3_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_evalue_weight: folded_blocks_0_stream_blocks_3_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_value_weight_valid: folded_blocks_0_stream_blocks_3_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_3_attention_value_bias_valid, folded_blocks_0_stream_blocks_3_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_3_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_3_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_mvalue_bias: folded_blocks_0_stream_blocks_3_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_evalue_bias: folded_blocks_0_stream_blocks_3_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_value_bias_valid: folded_blocks_0_stream_blocks_3_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_3_attention_proj_weight_valid, folded_blocks_0_stream_blocks_3_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_3_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_3_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_mproj_weight: folded_blocks_0_stream_blocks_3_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_eproj_weight: folded_blocks_0_stream_blocks_3_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_proj_weight_valid: folded_blocks_0_stream_blocks_3_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_3_attention_proj_bias_valid, folded_blocks_0_stream_blocks_3_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_3_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_3_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_mproj_bias: folded_blocks_0_stream_blocks_3_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_eproj_bias: folded_blocks_0_stream_blocks_3_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_attention_proj_bias_valid: folded_blocks_0_stream_blocks_3_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_norm2_eweight;
logic folded_blocks_0_stream_blocks_3_norm2_weight_valid, folded_blocks_0_stream_blocks_3_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_3_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_3_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm2_mweight: folded_blocks_0_stream_blocks_3_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm2_eweight: folded_blocks_0_stream_blocks_3_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm2_weight_valid: folded_blocks_0_stream_blocks_3_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_3_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_3_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_3_norm2_ebias;
logic folded_blocks_0_stream_blocks_3_norm2_bias_valid, folded_blocks_0_stream_blocks_3_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_3_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_3_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_3_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_3_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_3_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_3_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_3_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm2_mbias: folded_blocks_0_stream_blocks_3_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm2_ebias: folded_blocks_0_stream_blocks_3_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_3_norm2_bias_valid: folded_blocks_0_stream_blocks_3_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_linear1_eweight;
logic folded_blocks_0_stream_blocks_4_linear1_weight_valid, folded_blocks_0_stream_blocks_4_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_4_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_4_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear1_mweight: folded_blocks_0_stream_blocks_4_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear1_eweight: folded_blocks_0_stream_blocks_4_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear1_weight_valid: folded_blocks_0_stream_blocks_4_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_linear1_ebias;
logic folded_blocks_0_stream_blocks_4_linear1_bias_valid, folded_blocks_0_stream_blocks_4_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_4_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_4_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear1_mbias: folded_blocks_0_stream_blocks_4_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear1_ebias: folded_blocks_0_stream_blocks_4_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear1_bias_valid: folded_blocks_0_stream_blocks_4_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_linear2_eweight;
logic folded_blocks_0_stream_blocks_4_linear2_weight_valid, folded_blocks_0_stream_blocks_4_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_4_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_4_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear2_mweight: folded_blocks_0_stream_blocks_4_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear2_eweight: folded_blocks_0_stream_blocks_4_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear2_weight_valid: folded_blocks_0_stream_blocks_4_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_linear2_ebias;
logic folded_blocks_0_stream_blocks_4_linear2_bias_valid, folded_blocks_0_stream_blocks_4_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_4_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_4_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear2_mbias: folded_blocks_0_stream_blocks_4_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear2_ebias: folded_blocks_0_stream_blocks_4_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_linear2_bias_valid: folded_blocks_0_stream_blocks_4_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_norm1_eweight;
logic folded_blocks_0_stream_blocks_4_norm1_weight_valid, folded_blocks_0_stream_blocks_4_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_4_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_4_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm1_mweight: folded_blocks_0_stream_blocks_4_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm1_eweight: folded_blocks_0_stream_blocks_4_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm1_weight_valid: folded_blocks_0_stream_blocks_4_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_norm1_ebias;
logic folded_blocks_0_stream_blocks_4_norm1_bias_valid, folded_blocks_0_stream_blocks_4_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_4_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_4_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm1_mbias: folded_blocks_0_stream_blocks_4_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm1_ebias: folded_blocks_0_stream_blocks_4_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm1_bias_valid: folded_blocks_0_stream_blocks_4_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_attention_equery_weight;
logic folded_blocks_0_stream_blocks_4_attention_query_weight_valid, folded_blocks_0_stream_blocks_4_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_4_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_4_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_mquery_weight: folded_blocks_0_stream_blocks_4_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_equery_weight: folded_blocks_0_stream_blocks_4_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_query_weight_valid: folded_blocks_0_stream_blocks_4_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_attention_equery_bias;
logic folded_blocks_0_stream_blocks_4_attention_query_bias_valid, folded_blocks_0_stream_blocks_4_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_4_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_4_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_mquery_bias: folded_blocks_0_stream_blocks_4_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_equery_bias: folded_blocks_0_stream_blocks_4_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_query_bias_valid: folded_blocks_0_stream_blocks_4_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_4_attention_key_weight_valid, folded_blocks_0_stream_blocks_4_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_4_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_4_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_mkey_weight: folded_blocks_0_stream_blocks_4_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_ekey_weight: folded_blocks_0_stream_blocks_4_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_key_weight_valid: folded_blocks_0_stream_blocks_4_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_4_attention_key_bias_valid, folded_blocks_0_stream_blocks_4_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_4_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_4_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_mkey_bias: folded_blocks_0_stream_blocks_4_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_ekey_bias: folded_blocks_0_stream_blocks_4_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_key_bias_valid: folded_blocks_0_stream_blocks_4_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_4_attention_value_weight_valid, folded_blocks_0_stream_blocks_4_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_4_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_4_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_mvalue_weight: folded_blocks_0_stream_blocks_4_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_evalue_weight: folded_blocks_0_stream_blocks_4_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_value_weight_valid: folded_blocks_0_stream_blocks_4_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_4_attention_value_bias_valid, folded_blocks_0_stream_blocks_4_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_4_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_4_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_mvalue_bias: folded_blocks_0_stream_blocks_4_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_evalue_bias: folded_blocks_0_stream_blocks_4_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_value_bias_valid: folded_blocks_0_stream_blocks_4_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_4_attention_proj_weight_valid, folded_blocks_0_stream_blocks_4_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_4_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_4_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_mproj_weight: folded_blocks_0_stream_blocks_4_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_eproj_weight: folded_blocks_0_stream_blocks_4_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_proj_weight_valid: folded_blocks_0_stream_blocks_4_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_4_attention_proj_bias_valid, folded_blocks_0_stream_blocks_4_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_4_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_4_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_mproj_bias: folded_blocks_0_stream_blocks_4_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_eproj_bias: folded_blocks_0_stream_blocks_4_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_attention_proj_bias_valid: folded_blocks_0_stream_blocks_4_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_norm2_eweight;
logic folded_blocks_0_stream_blocks_4_norm2_weight_valid, folded_blocks_0_stream_blocks_4_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_4_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_4_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm2_mweight: folded_blocks_0_stream_blocks_4_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm2_eweight: folded_blocks_0_stream_blocks_4_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm2_weight_valid: folded_blocks_0_stream_blocks_4_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_4_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_4_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_4_norm2_ebias;
logic folded_blocks_0_stream_blocks_4_norm2_bias_valid, folded_blocks_0_stream_blocks_4_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_4_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_4_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_4_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_4_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_4_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_4_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_4_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm2_mbias: folded_blocks_0_stream_blocks_4_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm2_ebias: folded_blocks_0_stream_blocks_4_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_4_norm2_bias_valid: folded_blocks_0_stream_blocks_4_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_linear1_eweight;
logic folded_blocks_0_stream_blocks_5_linear1_weight_valid, folded_blocks_0_stream_blocks_5_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_5_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_5_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear1_mweight: folded_blocks_0_stream_blocks_5_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear1_eweight: folded_blocks_0_stream_blocks_5_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear1_weight_valid: folded_blocks_0_stream_blocks_5_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_linear1_ebias;
logic folded_blocks_0_stream_blocks_5_linear1_bias_valid, folded_blocks_0_stream_blocks_5_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_5_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_5_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear1_mbias: folded_blocks_0_stream_blocks_5_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear1_ebias: folded_blocks_0_stream_blocks_5_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear1_bias_valid: folded_blocks_0_stream_blocks_5_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_linear2_eweight;
logic folded_blocks_0_stream_blocks_5_linear2_weight_valid, folded_blocks_0_stream_blocks_5_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_5_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_5_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear2_mweight: folded_blocks_0_stream_blocks_5_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear2_eweight: folded_blocks_0_stream_blocks_5_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear2_weight_valid: folded_blocks_0_stream_blocks_5_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_linear2_ebias;
logic folded_blocks_0_stream_blocks_5_linear2_bias_valid, folded_blocks_0_stream_blocks_5_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_5_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_5_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear2_mbias: folded_blocks_0_stream_blocks_5_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear2_ebias: folded_blocks_0_stream_blocks_5_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_linear2_bias_valid: folded_blocks_0_stream_blocks_5_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_norm1_eweight;
logic folded_blocks_0_stream_blocks_5_norm1_weight_valid, folded_blocks_0_stream_blocks_5_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_5_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_5_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm1_mweight: folded_blocks_0_stream_blocks_5_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm1_eweight: folded_blocks_0_stream_blocks_5_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm1_weight_valid: folded_blocks_0_stream_blocks_5_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_norm1_ebias;
logic folded_blocks_0_stream_blocks_5_norm1_bias_valid, folded_blocks_0_stream_blocks_5_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_5_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_5_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm1_mbias: folded_blocks_0_stream_blocks_5_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm1_ebias: folded_blocks_0_stream_blocks_5_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm1_bias_valid: folded_blocks_0_stream_blocks_5_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_attention_equery_weight;
logic folded_blocks_0_stream_blocks_5_attention_query_weight_valid, folded_blocks_0_stream_blocks_5_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_5_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_5_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_mquery_weight: folded_blocks_0_stream_blocks_5_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_equery_weight: folded_blocks_0_stream_blocks_5_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_query_weight_valid: folded_blocks_0_stream_blocks_5_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_attention_equery_bias;
logic folded_blocks_0_stream_blocks_5_attention_query_bias_valid, folded_blocks_0_stream_blocks_5_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_5_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_5_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_mquery_bias: folded_blocks_0_stream_blocks_5_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_equery_bias: folded_blocks_0_stream_blocks_5_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_query_bias_valid: folded_blocks_0_stream_blocks_5_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_5_attention_key_weight_valid, folded_blocks_0_stream_blocks_5_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_5_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_5_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_mkey_weight: folded_blocks_0_stream_blocks_5_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_ekey_weight: folded_blocks_0_stream_blocks_5_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_key_weight_valid: folded_blocks_0_stream_blocks_5_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_5_attention_key_bias_valid, folded_blocks_0_stream_blocks_5_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_5_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_5_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_mkey_bias: folded_blocks_0_stream_blocks_5_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_ekey_bias: folded_blocks_0_stream_blocks_5_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_key_bias_valid: folded_blocks_0_stream_blocks_5_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_5_attention_value_weight_valid, folded_blocks_0_stream_blocks_5_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_5_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_5_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_mvalue_weight: folded_blocks_0_stream_blocks_5_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_evalue_weight: folded_blocks_0_stream_blocks_5_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_value_weight_valid: folded_blocks_0_stream_blocks_5_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_5_attention_value_bias_valid, folded_blocks_0_stream_blocks_5_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_5_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_5_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_mvalue_bias: folded_blocks_0_stream_blocks_5_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_evalue_bias: folded_blocks_0_stream_blocks_5_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_value_bias_valid: folded_blocks_0_stream_blocks_5_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_5_attention_proj_weight_valid, folded_blocks_0_stream_blocks_5_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_5_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_5_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_mproj_weight: folded_blocks_0_stream_blocks_5_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_eproj_weight: folded_blocks_0_stream_blocks_5_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_proj_weight_valid: folded_blocks_0_stream_blocks_5_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_5_attention_proj_bias_valid, folded_blocks_0_stream_blocks_5_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_5_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_5_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_mproj_bias: folded_blocks_0_stream_blocks_5_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_eproj_bias: folded_blocks_0_stream_blocks_5_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_attention_proj_bias_valid: folded_blocks_0_stream_blocks_5_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_norm2_eweight;
logic folded_blocks_0_stream_blocks_5_norm2_weight_valid, folded_blocks_0_stream_blocks_5_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_5_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_5_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm2_mweight: folded_blocks_0_stream_blocks_5_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm2_eweight: folded_blocks_0_stream_blocks_5_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm2_weight_valid: folded_blocks_0_stream_blocks_5_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_5_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_5_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_5_norm2_ebias;
logic folded_blocks_0_stream_blocks_5_norm2_bias_valid, folded_blocks_0_stream_blocks_5_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_5_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_5_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_5_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_5_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_5_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_5_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_5_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm2_mbias: folded_blocks_0_stream_blocks_5_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm2_ebias: folded_blocks_0_stream_blocks_5_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_5_norm2_bias_valid: folded_blocks_0_stream_blocks_5_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_linear1_eweight;
logic folded_blocks_0_stream_blocks_6_linear1_weight_valid, folded_blocks_0_stream_blocks_6_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_6_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_6_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear1_mweight: folded_blocks_0_stream_blocks_6_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear1_eweight: folded_blocks_0_stream_blocks_6_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear1_weight_valid: folded_blocks_0_stream_blocks_6_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_linear1_ebias;
logic folded_blocks_0_stream_blocks_6_linear1_bias_valid, folded_blocks_0_stream_blocks_6_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_6_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_6_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear1_mbias: folded_blocks_0_stream_blocks_6_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear1_ebias: folded_blocks_0_stream_blocks_6_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear1_bias_valid: folded_blocks_0_stream_blocks_6_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_linear2_eweight;
logic folded_blocks_0_stream_blocks_6_linear2_weight_valid, folded_blocks_0_stream_blocks_6_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_6_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_6_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear2_mweight: folded_blocks_0_stream_blocks_6_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear2_eweight: folded_blocks_0_stream_blocks_6_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear2_weight_valid: folded_blocks_0_stream_blocks_6_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_linear2_ebias;
logic folded_blocks_0_stream_blocks_6_linear2_bias_valid, folded_blocks_0_stream_blocks_6_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_6_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_6_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear2_mbias: folded_blocks_0_stream_blocks_6_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear2_ebias: folded_blocks_0_stream_blocks_6_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_linear2_bias_valid: folded_blocks_0_stream_blocks_6_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_norm1_eweight;
logic folded_blocks_0_stream_blocks_6_norm1_weight_valid, folded_blocks_0_stream_blocks_6_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_6_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_6_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm1_mweight: folded_blocks_0_stream_blocks_6_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm1_eweight: folded_blocks_0_stream_blocks_6_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm1_weight_valid: folded_blocks_0_stream_blocks_6_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_norm1_ebias;
logic folded_blocks_0_stream_blocks_6_norm1_bias_valid, folded_blocks_0_stream_blocks_6_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_6_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_6_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm1_mbias: folded_blocks_0_stream_blocks_6_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm1_ebias: folded_blocks_0_stream_blocks_6_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm1_bias_valid: folded_blocks_0_stream_blocks_6_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_attention_equery_weight;
logic folded_blocks_0_stream_blocks_6_attention_query_weight_valid, folded_blocks_0_stream_blocks_6_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_6_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_6_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_mquery_weight: folded_blocks_0_stream_blocks_6_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_equery_weight: folded_blocks_0_stream_blocks_6_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_query_weight_valid: folded_blocks_0_stream_blocks_6_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_attention_equery_bias;
logic folded_blocks_0_stream_blocks_6_attention_query_bias_valid, folded_blocks_0_stream_blocks_6_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_6_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_6_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_mquery_bias: folded_blocks_0_stream_blocks_6_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_equery_bias: folded_blocks_0_stream_blocks_6_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_query_bias_valid: folded_blocks_0_stream_blocks_6_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_6_attention_key_weight_valid, folded_blocks_0_stream_blocks_6_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_6_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_6_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_mkey_weight: folded_blocks_0_stream_blocks_6_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_ekey_weight: folded_blocks_0_stream_blocks_6_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_key_weight_valid: folded_blocks_0_stream_blocks_6_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_6_attention_key_bias_valid, folded_blocks_0_stream_blocks_6_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_6_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_6_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_mkey_bias: folded_blocks_0_stream_blocks_6_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_ekey_bias: folded_blocks_0_stream_blocks_6_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_key_bias_valid: folded_blocks_0_stream_blocks_6_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_6_attention_value_weight_valid, folded_blocks_0_stream_blocks_6_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_6_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_6_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_mvalue_weight: folded_blocks_0_stream_blocks_6_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_evalue_weight: folded_blocks_0_stream_blocks_6_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_value_weight_valid: folded_blocks_0_stream_blocks_6_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_6_attention_value_bias_valid, folded_blocks_0_stream_blocks_6_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_6_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_6_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_mvalue_bias: folded_blocks_0_stream_blocks_6_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_evalue_bias: folded_blocks_0_stream_blocks_6_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_value_bias_valid: folded_blocks_0_stream_blocks_6_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_6_attention_proj_weight_valid, folded_blocks_0_stream_blocks_6_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_6_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_6_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_mproj_weight: folded_blocks_0_stream_blocks_6_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_eproj_weight: folded_blocks_0_stream_blocks_6_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_proj_weight_valid: folded_blocks_0_stream_blocks_6_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_6_attention_proj_bias_valid, folded_blocks_0_stream_blocks_6_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_6_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_6_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_mproj_bias: folded_blocks_0_stream_blocks_6_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_eproj_bias: folded_blocks_0_stream_blocks_6_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_attention_proj_bias_valid: folded_blocks_0_stream_blocks_6_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_norm2_eweight;
logic folded_blocks_0_stream_blocks_6_norm2_weight_valid, folded_blocks_0_stream_blocks_6_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_6_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_6_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm2_mweight: folded_blocks_0_stream_blocks_6_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm2_eweight: folded_blocks_0_stream_blocks_6_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm2_weight_valid: folded_blocks_0_stream_blocks_6_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_6_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_6_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_6_norm2_ebias;
logic folded_blocks_0_stream_blocks_6_norm2_bias_valid, folded_blocks_0_stream_blocks_6_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_6_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_6_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_6_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_6_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_6_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_6_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_6_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm2_mbias: folded_blocks_0_stream_blocks_6_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm2_ebias: folded_blocks_0_stream_blocks_6_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_6_norm2_bias_valid: folded_blocks_0_stream_blocks_6_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_linear1_eweight;
logic folded_blocks_0_stream_blocks_7_linear1_weight_valid, folded_blocks_0_stream_blocks_7_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_7_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_7_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear1_mweight: folded_blocks_0_stream_blocks_7_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear1_eweight: folded_blocks_0_stream_blocks_7_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear1_weight_valid: folded_blocks_0_stream_blocks_7_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_linear1_ebias;
logic folded_blocks_0_stream_blocks_7_linear1_bias_valid, folded_blocks_0_stream_blocks_7_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_7_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_7_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear1_mbias: folded_blocks_0_stream_blocks_7_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear1_ebias: folded_blocks_0_stream_blocks_7_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear1_bias_valid: folded_blocks_0_stream_blocks_7_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_linear2_eweight;
logic folded_blocks_0_stream_blocks_7_linear2_weight_valid, folded_blocks_0_stream_blocks_7_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_7_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_7_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear2_mweight: folded_blocks_0_stream_blocks_7_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear2_eweight: folded_blocks_0_stream_blocks_7_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear2_weight_valid: folded_blocks_0_stream_blocks_7_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_linear2_ebias;
logic folded_blocks_0_stream_blocks_7_linear2_bias_valid, folded_blocks_0_stream_blocks_7_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_7_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_7_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear2_mbias: folded_blocks_0_stream_blocks_7_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear2_ebias: folded_blocks_0_stream_blocks_7_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_linear2_bias_valid: folded_blocks_0_stream_blocks_7_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_norm1_eweight;
logic folded_blocks_0_stream_blocks_7_norm1_weight_valid, folded_blocks_0_stream_blocks_7_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_7_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_7_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm1_mweight: folded_blocks_0_stream_blocks_7_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm1_eweight: folded_blocks_0_stream_blocks_7_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm1_weight_valid: folded_blocks_0_stream_blocks_7_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_norm1_ebias;
logic folded_blocks_0_stream_blocks_7_norm1_bias_valid, folded_blocks_0_stream_blocks_7_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_7_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_7_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm1_mbias: folded_blocks_0_stream_blocks_7_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm1_ebias: folded_blocks_0_stream_blocks_7_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm1_bias_valid: folded_blocks_0_stream_blocks_7_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_attention_equery_weight;
logic folded_blocks_0_stream_blocks_7_attention_query_weight_valid, folded_blocks_0_stream_blocks_7_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_7_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_7_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_mquery_weight: folded_blocks_0_stream_blocks_7_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_equery_weight: folded_blocks_0_stream_blocks_7_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_query_weight_valid: folded_blocks_0_stream_blocks_7_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_attention_equery_bias;
logic folded_blocks_0_stream_blocks_7_attention_query_bias_valid, folded_blocks_0_stream_blocks_7_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_7_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_7_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_mquery_bias: folded_blocks_0_stream_blocks_7_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_equery_bias: folded_blocks_0_stream_blocks_7_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_query_bias_valid: folded_blocks_0_stream_blocks_7_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_7_attention_key_weight_valid, folded_blocks_0_stream_blocks_7_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_7_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_7_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_mkey_weight: folded_blocks_0_stream_blocks_7_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_ekey_weight: folded_blocks_0_stream_blocks_7_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_key_weight_valid: folded_blocks_0_stream_blocks_7_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_7_attention_key_bias_valid, folded_blocks_0_stream_blocks_7_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_7_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_7_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_mkey_bias: folded_blocks_0_stream_blocks_7_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_ekey_bias: folded_blocks_0_stream_blocks_7_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_key_bias_valid: folded_blocks_0_stream_blocks_7_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_7_attention_value_weight_valid, folded_blocks_0_stream_blocks_7_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_7_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_7_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_mvalue_weight: folded_blocks_0_stream_blocks_7_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_evalue_weight: folded_blocks_0_stream_blocks_7_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_value_weight_valid: folded_blocks_0_stream_blocks_7_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_7_attention_value_bias_valid, folded_blocks_0_stream_blocks_7_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_7_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_7_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_mvalue_bias: folded_blocks_0_stream_blocks_7_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_evalue_bias: folded_blocks_0_stream_blocks_7_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_value_bias_valid: folded_blocks_0_stream_blocks_7_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_7_attention_proj_weight_valid, folded_blocks_0_stream_blocks_7_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_7_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_7_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_mproj_weight: folded_blocks_0_stream_blocks_7_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_eproj_weight: folded_blocks_0_stream_blocks_7_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_proj_weight_valid: folded_blocks_0_stream_blocks_7_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_7_attention_proj_bias_valid, folded_blocks_0_stream_blocks_7_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_7_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_7_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_mproj_bias: folded_blocks_0_stream_blocks_7_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_eproj_bias: folded_blocks_0_stream_blocks_7_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_attention_proj_bias_valid: folded_blocks_0_stream_blocks_7_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_norm2_eweight;
logic folded_blocks_0_stream_blocks_7_norm2_weight_valid, folded_blocks_0_stream_blocks_7_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_7_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_7_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm2_mweight: folded_blocks_0_stream_blocks_7_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm2_eweight: folded_blocks_0_stream_blocks_7_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm2_weight_valid: folded_blocks_0_stream_blocks_7_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_7_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_7_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_7_norm2_ebias;
logic folded_blocks_0_stream_blocks_7_norm2_bias_valid, folded_blocks_0_stream_blocks_7_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_7_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_7_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_7_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_7_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_7_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_7_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_7_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm2_mbias: folded_blocks_0_stream_blocks_7_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm2_ebias: folded_blocks_0_stream_blocks_7_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_7_norm2_bias_valid: folded_blocks_0_stream_blocks_7_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_linear1_eweight;
logic folded_blocks_0_stream_blocks_8_linear1_weight_valid, folded_blocks_0_stream_blocks_8_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_8_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_8_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear1_mweight: folded_blocks_0_stream_blocks_8_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear1_eweight: folded_blocks_0_stream_blocks_8_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear1_weight_valid: folded_blocks_0_stream_blocks_8_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_linear1_ebias;
logic folded_blocks_0_stream_blocks_8_linear1_bias_valid, folded_blocks_0_stream_blocks_8_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_8_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_8_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear1_mbias: folded_blocks_0_stream_blocks_8_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear1_ebias: folded_blocks_0_stream_blocks_8_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear1_bias_valid: folded_blocks_0_stream_blocks_8_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_linear2_eweight;
logic folded_blocks_0_stream_blocks_8_linear2_weight_valid, folded_blocks_0_stream_blocks_8_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_8_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_8_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear2_mweight: folded_blocks_0_stream_blocks_8_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear2_eweight: folded_blocks_0_stream_blocks_8_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear2_weight_valid: folded_blocks_0_stream_blocks_8_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_linear2_ebias;
logic folded_blocks_0_stream_blocks_8_linear2_bias_valid, folded_blocks_0_stream_blocks_8_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_8_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_8_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear2_mbias: folded_blocks_0_stream_blocks_8_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear2_ebias: folded_blocks_0_stream_blocks_8_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_linear2_bias_valid: folded_blocks_0_stream_blocks_8_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_norm1_eweight;
logic folded_blocks_0_stream_blocks_8_norm1_weight_valid, folded_blocks_0_stream_blocks_8_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_8_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_8_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm1_mweight: folded_blocks_0_stream_blocks_8_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm1_eweight: folded_blocks_0_stream_blocks_8_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm1_weight_valid: folded_blocks_0_stream_blocks_8_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_norm1_ebias;
logic folded_blocks_0_stream_blocks_8_norm1_bias_valid, folded_blocks_0_stream_blocks_8_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_8_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_8_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm1_mbias: folded_blocks_0_stream_blocks_8_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm1_ebias: folded_blocks_0_stream_blocks_8_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm1_bias_valid: folded_blocks_0_stream_blocks_8_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_attention_equery_weight;
logic folded_blocks_0_stream_blocks_8_attention_query_weight_valid, folded_blocks_0_stream_blocks_8_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_8_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_8_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_mquery_weight: folded_blocks_0_stream_blocks_8_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_equery_weight: folded_blocks_0_stream_blocks_8_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_query_weight_valid: folded_blocks_0_stream_blocks_8_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_attention_equery_bias;
logic folded_blocks_0_stream_blocks_8_attention_query_bias_valid, folded_blocks_0_stream_blocks_8_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_8_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_8_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_mquery_bias: folded_blocks_0_stream_blocks_8_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_equery_bias: folded_blocks_0_stream_blocks_8_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_query_bias_valid: folded_blocks_0_stream_blocks_8_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_8_attention_key_weight_valid, folded_blocks_0_stream_blocks_8_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_8_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_8_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_mkey_weight: folded_blocks_0_stream_blocks_8_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_ekey_weight: folded_blocks_0_stream_blocks_8_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_key_weight_valid: folded_blocks_0_stream_blocks_8_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_8_attention_key_bias_valid, folded_blocks_0_stream_blocks_8_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_8_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_8_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_mkey_bias: folded_blocks_0_stream_blocks_8_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_ekey_bias: folded_blocks_0_stream_blocks_8_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_key_bias_valid: folded_blocks_0_stream_blocks_8_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_8_attention_value_weight_valid, folded_blocks_0_stream_blocks_8_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_8_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_8_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_mvalue_weight: folded_blocks_0_stream_blocks_8_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_evalue_weight: folded_blocks_0_stream_blocks_8_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_value_weight_valid: folded_blocks_0_stream_blocks_8_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_8_attention_value_bias_valid, folded_blocks_0_stream_blocks_8_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_8_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_8_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_mvalue_bias: folded_blocks_0_stream_blocks_8_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_evalue_bias: folded_blocks_0_stream_blocks_8_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_value_bias_valid: folded_blocks_0_stream_blocks_8_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_8_attention_proj_weight_valid, folded_blocks_0_stream_blocks_8_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_8_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_8_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_mproj_weight: folded_blocks_0_stream_blocks_8_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_eproj_weight: folded_blocks_0_stream_blocks_8_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_proj_weight_valid: folded_blocks_0_stream_blocks_8_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_8_attention_proj_bias_valid, folded_blocks_0_stream_blocks_8_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_8_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_8_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_mproj_bias: folded_blocks_0_stream_blocks_8_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_eproj_bias: folded_blocks_0_stream_blocks_8_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_attention_proj_bias_valid: folded_blocks_0_stream_blocks_8_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_norm2_eweight;
logic folded_blocks_0_stream_blocks_8_norm2_weight_valid, folded_blocks_0_stream_blocks_8_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_8_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_8_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm2_mweight: folded_blocks_0_stream_blocks_8_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm2_eweight: folded_blocks_0_stream_blocks_8_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm2_weight_valid: folded_blocks_0_stream_blocks_8_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_8_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_8_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_8_norm2_ebias;
logic folded_blocks_0_stream_blocks_8_norm2_bias_valid, folded_blocks_0_stream_blocks_8_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_8_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_8_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_8_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_8_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_8_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_8_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_8_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm2_mbias: folded_blocks_0_stream_blocks_8_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm2_ebias: folded_blocks_0_stream_blocks_8_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_8_norm2_bias_valid: folded_blocks_0_stream_blocks_8_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_linear1_eweight;
logic folded_blocks_0_stream_blocks_9_linear1_weight_valid, folded_blocks_0_stream_blocks_9_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_9_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_9_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear1_mweight: folded_blocks_0_stream_blocks_9_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear1_eweight: folded_blocks_0_stream_blocks_9_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear1_weight_valid: folded_blocks_0_stream_blocks_9_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_linear1_ebias;
logic folded_blocks_0_stream_blocks_9_linear1_bias_valid, folded_blocks_0_stream_blocks_9_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_9_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_9_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear1_mbias: folded_blocks_0_stream_blocks_9_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear1_ebias: folded_blocks_0_stream_blocks_9_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear1_bias_valid: folded_blocks_0_stream_blocks_9_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_linear2_eweight;
logic folded_blocks_0_stream_blocks_9_linear2_weight_valid, folded_blocks_0_stream_blocks_9_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_9_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_9_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear2_mweight: folded_blocks_0_stream_blocks_9_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear2_eweight: folded_blocks_0_stream_blocks_9_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear2_weight_valid: folded_blocks_0_stream_blocks_9_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_linear2_ebias;
logic folded_blocks_0_stream_blocks_9_linear2_bias_valid, folded_blocks_0_stream_blocks_9_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_9_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_9_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear2_mbias: folded_blocks_0_stream_blocks_9_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear2_ebias: folded_blocks_0_stream_blocks_9_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_linear2_bias_valid: folded_blocks_0_stream_blocks_9_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_norm1_eweight;
logic folded_blocks_0_stream_blocks_9_norm1_weight_valid, folded_blocks_0_stream_blocks_9_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_9_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_9_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm1_mweight: folded_blocks_0_stream_blocks_9_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm1_eweight: folded_blocks_0_stream_blocks_9_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm1_weight_valid: folded_blocks_0_stream_blocks_9_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_norm1_ebias;
logic folded_blocks_0_stream_blocks_9_norm1_bias_valid, folded_blocks_0_stream_blocks_9_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_9_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_9_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm1_mbias: folded_blocks_0_stream_blocks_9_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm1_ebias: folded_blocks_0_stream_blocks_9_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm1_bias_valid: folded_blocks_0_stream_blocks_9_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_attention_equery_weight;
logic folded_blocks_0_stream_blocks_9_attention_query_weight_valid, folded_blocks_0_stream_blocks_9_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_9_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_9_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_mquery_weight: folded_blocks_0_stream_blocks_9_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_equery_weight: folded_blocks_0_stream_blocks_9_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_query_weight_valid: folded_blocks_0_stream_blocks_9_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_attention_equery_bias;
logic folded_blocks_0_stream_blocks_9_attention_query_bias_valid, folded_blocks_0_stream_blocks_9_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_9_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_9_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_mquery_bias: folded_blocks_0_stream_blocks_9_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_equery_bias: folded_blocks_0_stream_blocks_9_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_query_bias_valid: folded_blocks_0_stream_blocks_9_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_9_attention_key_weight_valid, folded_blocks_0_stream_blocks_9_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_9_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_9_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_mkey_weight: folded_blocks_0_stream_blocks_9_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_ekey_weight: folded_blocks_0_stream_blocks_9_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_key_weight_valid: folded_blocks_0_stream_blocks_9_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_9_attention_key_bias_valid, folded_blocks_0_stream_blocks_9_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_9_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_9_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_mkey_bias: folded_blocks_0_stream_blocks_9_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_ekey_bias: folded_blocks_0_stream_blocks_9_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_key_bias_valid: folded_blocks_0_stream_blocks_9_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_9_attention_value_weight_valid, folded_blocks_0_stream_blocks_9_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_9_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_9_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_mvalue_weight: folded_blocks_0_stream_blocks_9_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_evalue_weight: folded_blocks_0_stream_blocks_9_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_value_weight_valid: folded_blocks_0_stream_blocks_9_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_9_attention_value_bias_valid, folded_blocks_0_stream_blocks_9_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_9_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_9_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_mvalue_bias: folded_blocks_0_stream_blocks_9_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_evalue_bias: folded_blocks_0_stream_blocks_9_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_value_bias_valid: folded_blocks_0_stream_blocks_9_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_9_attention_proj_weight_valid, folded_blocks_0_stream_blocks_9_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_9_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_9_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_mproj_weight: folded_blocks_0_stream_blocks_9_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_eproj_weight: folded_blocks_0_stream_blocks_9_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_proj_weight_valid: folded_blocks_0_stream_blocks_9_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_9_attention_proj_bias_valid, folded_blocks_0_stream_blocks_9_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_9_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_9_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_mproj_bias: folded_blocks_0_stream_blocks_9_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_eproj_bias: folded_blocks_0_stream_blocks_9_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_attention_proj_bias_valid: folded_blocks_0_stream_blocks_9_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_norm2_eweight;
logic folded_blocks_0_stream_blocks_9_norm2_weight_valid, folded_blocks_0_stream_blocks_9_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_9_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_9_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm2_mweight: folded_blocks_0_stream_blocks_9_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm2_eweight: folded_blocks_0_stream_blocks_9_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm2_weight_valid: folded_blocks_0_stream_blocks_9_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_9_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_9_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_9_norm2_ebias;
logic folded_blocks_0_stream_blocks_9_norm2_bias_valid, folded_blocks_0_stream_blocks_9_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_9_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_9_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_9_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_9_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_9_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_9_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_9_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm2_mbias: folded_blocks_0_stream_blocks_9_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm2_ebias: folded_blocks_0_stream_blocks_9_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_9_norm2_bias_valid: folded_blocks_0_stream_blocks_9_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_linear1_eweight;
logic folded_blocks_0_stream_blocks_10_linear1_weight_valid, folded_blocks_0_stream_blocks_10_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_10_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_10_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear1_mweight: folded_blocks_0_stream_blocks_10_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear1_eweight: folded_blocks_0_stream_blocks_10_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear1_weight_valid: folded_blocks_0_stream_blocks_10_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_linear1_ebias;
logic folded_blocks_0_stream_blocks_10_linear1_bias_valid, folded_blocks_0_stream_blocks_10_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_10_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_10_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear1_mbias: folded_blocks_0_stream_blocks_10_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear1_ebias: folded_blocks_0_stream_blocks_10_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear1_bias_valid: folded_blocks_0_stream_blocks_10_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_linear2_eweight;
logic folded_blocks_0_stream_blocks_10_linear2_weight_valid, folded_blocks_0_stream_blocks_10_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_10_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_10_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear2_mweight: folded_blocks_0_stream_blocks_10_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear2_eweight: folded_blocks_0_stream_blocks_10_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear2_weight_valid: folded_blocks_0_stream_blocks_10_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_linear2_ebias;
logic folded_blocks_0_stream_blocks_10_linear2_bias_valid, folded_blocks_0_stream_blocks_10_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_10_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_10_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear2_mbias: folded_blocks_0_stream_blocks_10_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear2_ebias: folded_blocks_0_stream_blocks_10_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_linear2_bias_valid: folded_blocks_0_stream_blocks_10_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_norm1_eweight;
logic folded_blocks_0_stream_blocks_10_norm1_weight_valid, folded_blocks_0_stream_blocks_10_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_10_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_10_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm1_mweight: folded_blocks_0_stream_blocks_10_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm1_eweight: folded_blocks_0_stream_blocks_10_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm1_weight_valid: folded_blocks_0_stream_blocks_10_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_norm1_ebias;
logic folded_blocks_0_stream_blocks_10_norm1_bias_valid, folded_blocks_0_stream_blocks_10_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_10_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_10_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm1_mbias: folded_blocks_0_stream_blocks_10_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm1_ebias: folded_blocks_0_stream_blocks_10_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm1_bias_valid: folded_blocks_0_stream_blocks_10_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_attention_equery_weight;
logic folded_blocks_0_stream_blocks_10_attention_query_weight_valid, folded_blocks_0_stream_blocks_10_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_10_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_10_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_mquery_weight: folded_blocks_0_stream_blocks_10_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_equery_weight: folded_blocks_0_stream_blocks_10_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_query_weight_valid: folded_blocks_0_stream_blocks_10_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_attention_equery_bias;
logic folded_blocks_0_stream_blocks_10_attention_query_bias_valid, folded_blocks_0_stream_blocks_10_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_10_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_10_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_mquery_bias: folded_blocks_0_stream_blocks_10_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_equery_bias: folded_blocks_0_stream_blocks_10_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_query_bias_valid: folded_blocks_0_stream_blocks_10_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_10_attention_key_weight_valid, folded_blocks_0_stream_blocks_10_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_10_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_10_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_mkey_weight: folded_blocks_0_stream_blocks_10_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_ekey_weight: folded_blocks_0_stream_blocks_10_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_key_weight_valid: folded_blocks_0_stream_blocks_10_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_10_attention_key_bias_valid, folded_blocks_0_stream_blocks_10_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_10_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_10_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_mkey_bias: folded_blocks_0_stream_blocks_10_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_ekey_bias: folded_blocks_0_stream_blocks_10_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_key_bias_valid: folded_blocks_0_stream_blocks_10_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_10_attention_value_weight_valid, folded_blocks_0_stream_blocks_10_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_10_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_10_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_mvalue_weight: folded_blocks_0_stream_blocks_10_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_evalue_weight: folded_blocks_0_stream_blocks_10_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_value_weight_valid: folded_blocks_0_stream_blocks_10_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_10_attention_value_bias_valid, folded_blocks_0_stream_blocks_10_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_10_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_10_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_mvalue_bias: folded_blocks_0_stream_blocks_10_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_evalue_bias: folded_blocks_0_stream_blocks_10_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_value_bias_valid: folded_blocks_0_stream_blocks_10_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_10_attention_proj_weight_valid, folded_blocks_0_stream_blocks_10_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_10_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_10_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_mproj_weight: folded_blocks_0_stream_blocks_10_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_eproj_weight: folded_blocks_0_stream_blocks_10_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_proj_weight_valid: folded_blocks_0_stream_blocks_10_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_10_attention_proj_bias_valid, folded_blocks_0_stream_blocks_10_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_10_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_10_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_mproj_bias: folded_blocks_0_stream_blocks_10_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_eproj_bias: folded_blocks_0_stream_blocks_10_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_attention_proj_bias_valid: folded_blocks_0_stream_blocks_10_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_norm2_eweight;
logic folded_blocks_0_stream_blocks_10_norm2_weight_valid, folded_blocks_0_stream_blocks_10_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_10_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_10_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm2_mweight: folded_blocks_0_stream_blocks_10_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm2_eweight: folded_blocks_0_stream_blocks_10_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm2_weight_valid: folded_blocks_0_stream_blocks_10_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_10_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_10_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_10_norm2_ebias;
logic folded_blocks_0_stream_blocks_10_norm2_bias_valid, folded_blocks_0_stream_blocks_10_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_10_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_10_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_10_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_10_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_10_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_10_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_10_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm2_mbias: folded_blocks_0_stream_blocks_10_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm2_ebias: folded_blocks_0_stream_blocks_10_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_10_norm2_bias_valid: folded_blocks_0_stream_blocks_10_norm2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_linear1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_linear1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_linear1_eweight;
logic folded_blocks_0_stream_blocks_11_linear1_weight_valid, folded_blocks_0_stream_blocks_11_linear1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_linear1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_linear1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_linear1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_11_linear1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_11_linear1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_linear1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_linear1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear1_mweight: folded_blocks_0_stream_blocks_11_linear1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear1_eweight: folded_blocks_0_stream_blocks_11_linear1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear1_weight_valid: folded_blocks_0_stream_blocks_11_linear1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_linear1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 192;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_linear1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_linear1_ebias;
logic folded_blocks_0_stream_blocks_11_linear1_bias_valid, folded_blocks_0_stream_blocks_11_linear1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_linear1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_linear1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_linear1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_11_linear1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_11_linear1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_linear1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_linear1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear1_mbias: folded_blocks_0_stream_blocks_11_linear1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear1_ebias: folded_blocks_0_stream_blocks_11_linear1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear1_bias_valid: folded_blocks_0_stream_blocks_11_linear1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_linear2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 9216;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_linear2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_linear2_eweight;
logic folded_blocks_0_stream_blocks_11_linear2_weight_valid, folded_blocks_0_stream_blocks_11_linear2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_linear2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_linear2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_linear2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_11_linear2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_11_linear2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_linear2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_linear2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear2_mweight: folded_blocks_0_stream_blocks_11_linear2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear2_eweight: folded_blocks_0_stream_blocks_11_linear2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear2_weight_valid: folded_blocks_0_stream_blocks_11_linear2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_linear2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_linear2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_linear2_ebias;
logic folded_blocks_0_stream_blocks_11_linear2_bias_valid, folded_blocks_0_stream_blocks_11_linear2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_linear2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_linear2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_linear2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_11_linear2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_11_linear2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_linear2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_linear2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear2_mbias: folded_blocks_0_stream_blocks_11_linear2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear2_ebias: folded_blocks_0_stream_blocks_11_linear2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_linear2_bias_valid: folded_blocks_0_stream_blocks_11_linear2_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_norm1_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_norm1_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_norm1_eweight;
logic folded_blocks_0_stream_blocks_11_norm1_weight_valid, folded_blocks_0_stream_blocks_11_norm1_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_norm1_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_norm1_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_norm1_mweight),
    .edata_out(folded_blocks_0_stream_blocks_11_norm1_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_11_norm1_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_norm1_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_norm1_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm1_mweight: folded_blocks_0_stream_blocks_11_norm1_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm1_eweight: folded_blocks_0_stream_blocks_11_norm1_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm1_weight_valid: folded_blocks_0_stream_blocks_11_norm1_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_norm1_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_norm1_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_norm1_ebias;
logic folded_blocks_0_stream_blocks_11_norm1_bias_valid, folded_blocks_0_stream_blocks_11_norm1_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_norm1_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_norm1_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_norm1_mbias),
    .edata_out(folded_blocks_0_stream_blocks_11_norm1_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_11_norm1_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_norm1_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_norm1_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm1_mbias: folded_blocks_0_stream_blocks_11_norm1_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm1_ebias: folded_blocks_0_stream_blocks_11_norm1_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm1_bias_valid: folded_blocks_0_stream_blocks_11_norm1_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_attention_query_weight_source #(
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_WEIGHT_PRECISION_0 = -1,
    parameter QUERY_WEIGHT_PRECISION_1 = -1,

    parameter QUERY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter QUERY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_WEIGHT_PRECISION_0-1:0] mdata_out      [QUERY_WEIGHT_PARALLELISM_DIM_0 * QUERY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_attention_mquery_weight [QUERY_WEIGHT_PARALLELISM_DIM_0*QUERY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_attention_equery_weight;
logic folded_blocks_0_stream_blocks_11_attention_query_weight_valid, folded_blocks_0_stream_blocks_11_attention_query_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_attention_query_weight_source #(
    .QUERY_WEIGHT_PRECISION_0(QUERY_WEIGHT_PRECISION_0),
    .QUERY_WEIGHT_PRECISION_1(QUERY_WEIGHT_PRECISION_1),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_0(QUERY_WEIGHT_TENSOR_SIZE_DIM_0),
    .QUERY_WEIGHT_PARALLELISM_DIM_0(QUERY_WEIGHT_PARALLELISM_DIM_0),
    .QUERY_WEIGHT_TENSOR_SIZE_DIM_1(QUERY_WEIGHT_TENSOR_SIZE_DIM_1),
    .QUERY_WEIGHT_PARALLELISM_DIM_1(QUERY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_attention_query_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_attention_mquery_weight),
    .edata_out(folded_blocks_0_stream_blocks_11_attention_equery_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_11_attention_query_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_attention_query_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_attention_query_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_mquery_weight: folded_blocks_0_stream_blocks_11_attention_mquery_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_equery_weight: folded_blocks_0_stream_blocks_11_attention_equery_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_query_weight_valid: folded_blocks_0_stream_blocks_11_attention_query_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_attention_query_bias_source #(
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter QUERY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter QUERY_BIAS_PRECISION_0 = -1,
    parameter QUERY_BIAS_PRECISION_1 = -1,

    parameter QUERY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter QUERY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [QUERY_BIAS_PRECISION_0-1:0] mdata_out      [QUERY_BIAS_PARALLELISM_DIM_0 * QUERY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [QUERY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [QUERY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_attention_mquery_bias [QUERY_BIAS_PARALLELISM_DIM_0*QUERY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [QUERY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_attention_equery_bias;
logic folded_blocks_0_stream_blocks_11_attention_query_bias_valid, folded_blocks_0_stream_blocks_11_attention_query_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_attention_query_bias_source #(
    .QUERY_BIAS_PRECISION_0(QUERY_BIAS_PRECISION_0),
    .QUERY_BIAS_PRECISION_1(QUERY_BIAS_PRECISION_1),
    .QUERY_BIAS_TENSOR_SIZE_DIM_0(QUERY_BIAS_TENSOR_SIZE_DIM_0),
    .QUERY_BIAS_PARALLELISM_DIM_0(QUERY_BIAS_PARALLELISM_DIM_0),
    .QUERY_BIAS_TENSOR_SIZE_DIM_1(QUERY_BIAS_TENSOR_SIZE_DIM_1),
    .QUERY_BIAS_PARALLELISM_DIM_1(QUERY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_attention_query_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_attention_mquery_bias),
    .edata_out(folded_blocks_0_stream_blocks_11_attention_equery_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_11_attention_query_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_attention_query_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_attention_query_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_mquery_bias: folded_blocks_0_stream_blocks_11_attention_mquery_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_equery_bias: folded_blocks_0_stream_blocks_11_attention_equery_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_query_bias_valid: folded_blocks_0_stream_blocks_11_attention_query_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_attention_key_weight_source #(
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_WEIGHT_PRECISION_0 = -1,
    parameter KEY_WEIGHT_PRECISION_1 = -1,

    parameter KEY_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter KEY_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_WEIGHT_PRECISION_0-1:0] mdata_out      [KEY_WEIGHT_PARALLELISM_DIM_0 * KEY_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [KEY_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_attention_mkey_weight [KEY_WEIGHT_PARALLELISM_DIM_0*KEY_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [KEY_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_attention_ekey_weight;
logic folded_blocks_0_stream_blocks_11_attention_key_weight_valid, folded_blocks_0_stream_blocks_11_attention_key_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_attention_key_weight_source #(
    .KEY_WEIGHT_PRECISION_0(KEY_WEIGHT_PRECISION_0),
    .KEY_WEIGHT_PRECISION_1(KEY_WEIGHT_PRECISION_1),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_0(KEY_WEIGHT_TENSOR_SIZE_DIM_0),
    .KEY_WEIGHT_PARALLELISM_DIM_0(KEY_WEIGHT_PARALLELISM_DIM_0),
    .KEY_WEIGHT_TENSOR_SIZE_DIM_1(KEY_WEIGHT_TENSOR_SIZE_DIM_1),
    .KEY_WEIGHT_PARALLELISM_DIM_1(KEY_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_attention_key_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_attention_mkey_weight),
    .edata_out(folded_blocks_0_stream_blocks_11_attention_ekey_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_11_attention_key_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_attention_key_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_attention_key_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_mkey_weight: folded_blocks_0_stream_blocks_11_attention_mkey_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_ekey_weight: folded_blocks_0_stream_blocks_11_attention_ekey_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_key_weight_valid: folded_blocks_0_stream_blocks_11_attention_key_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_attention_key_bias_source #(
    parameter KEY_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter KEY_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter KEY_BIAS_PRECISION_0 = -1,
    parameter KEY_BIAS_PRECISION_1 = -1,

    parameter KEY_BIAS_PARALLELISM_DIM_0 = -1,
    parameter KEY_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [KEY_BIAS_PRECISION_0-1:0] mdata_out      [KEY_BIAS_PARALLELISM_DIM_0 * KEY_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [KEY_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [KEY_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_attention_mkey_bias [KEY_BIAS_PARALLELISM_DIM_0*KEY_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [KEY_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_attention_ekey_bias;
logic folded_blocks_0_stream_blocks_11_attention_key_bias_valid, folded_blocks_0_stream_blocks_11_attention_key_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_attention_key_bias_source #(
    .KEY_BIAS_PRECISION_0(KEY_BIAS_PRECISION_0),
    .KEY_BIAS_PRECISION_1(KEY_BIAS_PRECISION_1),
    .KEY_BIAS_TENSOR_SIZE_DIM_0(KEY_BIAS_TENSOR_SIZE_DIM_0),
    .KEY_BIAS_PARALLELISM_DIM_0(KEY_BIAS_PARALLELISM_DIM_0),
    .KEY_BIAS_TENSOR_SIZE_DIM_1(KEY_BIAS_TENSOR_SIZE_DIM_1),
    .KEY_BIAS_PARALLELISM_DIM_1(KEY_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_attention_key_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_attention_mkey_bias),
    .edata_out(folded_blocks_0_stream_blocks_11_attention_ekey_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_11_attention_key_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_attention_key_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_attention_key_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_mkey_bias: folded_blocks_0_stream_blocks_11_attention_mkey_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_ekey_bias: folded_blocks_0_stream_blocks_11_attention_ekey_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_key_bias_valid: folded_blocks_0_stream_blocks_11_attention_key_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_attention_value_weight_source #(
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_WEIGHT_PRECISION_0 = -1,
    parameter VALUE_WEIGHT_PRECISION_1 = -1,

    parameter VALUE_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter VALUE_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_WEIGHT_PRECISION_0-1:0] mdata_out      [VALUE_WEIGHT_PARALLELISM_DIM_0 * VALUE_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_attention_mvalue_weight [VALUE_WEIGHT_PARALLELISM_DIM_0*VALUE_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_attention_evalue_weight;
logic folded_blocks_0_stream_blocks_11_attention_value_weight_valid, folded_blocks_0_stream_blocks_11_attention_value_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_attention_value_weight_source #(
    .VALUE_WEIGHT_PRECISION_0(VALUE_WEIGHT_PRECISION_0),
    .VALUE_WEIGHT_PRECISION_1(VALUE_WEIGHT_PRECISION_1),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_0(VALUE_WEIGHT_TENSOR_SIZE_DIM_0),
    .VALUE_WEIGHT_PARALLELISM_DIM_0(VALUE_WEIGHT_PARALLELISM_DIM_0),
    .VALUE_WEIGHT_TENSOR_SIZE_DIM_1(VALUE_WEIGHT_TENSOR_SIZE_DIM_1),
    .VALUE_WEIGHT_PARALLELISM_DIM_1(VALUE_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_attention_value_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_attention_mvalue_weight),
    .edata_out(folded_blocks_0_stream_blocks_11_attention_evalue_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_11_attention_value_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_attention_value_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_attention_value_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_mvalue_weight: folded_blocks_0_stream_blocks_11_attention_mvalue_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_evalue_weight: folded_blocks_0_stream_blocks_11_attention_evalue_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_value_weight_valid: folded_blocks_0_stream_blocks_11_attention_value_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_attention_value_bias_source #(
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter VALUE_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter VALUE_BIAS_PRECISION_0 = -1,
    parameter VALUE_BIAS_PRECISION_1 = -1,

    parameter VALUE_BIAS_PARALLELISM_DIM_0 = -1,
    parameter VALUE_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [VALUE_BIAS_PRECISION_0-1:0] mdata_out      [VALUE_BIAS_PARALLELISM_DIM_0 * VALUE_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [VALUE_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [VALUE_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_attention_mvalue_bias [VALUE_BIAS_PARALLELISM_DIM_0*VALUE_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [VALUE_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_attention_evalue_bias;
logic folded_blocks_0_stream_blocks_11_attention_value_bias_valid, folded_blocks_0_stream_blocks_11_attention_value_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_attention_value_bias_source #(
    .VALUE_BIAS_PRECISION_0(VALUE_BIAS_PRECISION_0),
    .VALUE_BIAS_PRECISION_1(VALUE_BIAS_PRECISION_1),
    .VALUE_BIAS_TENSOR_SIZE_DIM_0(VALUE_BIAS_TENSOR_SIZE_DIM_0),
    .VALUE_BIAS_PARALLELISM_DIM_0(VALUE_BIAS_PARALLELISM_DIM_0),
    .VALUE_BIAS_TENSOR_SIZE_DIM_1(VALUE_BIAS_TENSOR_SIZE_DIM_1),
    .VALUE_BIAS_PARALLELISM_DIM_1(VALUE_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_attention_value_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_attention_mvalue_bias),
    .edata_out(folded_blocks_0_stream_blocks_11_attention_evalue_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_11_attention_value_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_attention_value_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_attention_value_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_mvalue_bias: folded_blocks_0_stream_blocks_11_attention_mvalue_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_evalue_bias: folded_blocks_0_stream_blocks_11_attention_evalue_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_value_bias_valid: folded_blocks_0_stream_blocks_11_attention_value_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_attention_proj_weight_source #(
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_WEIGHT_PRECISION_0 = -1,
    parameter PROJ_WEIGHT_PRECISION_1 = -1,

    parameter PROJ_WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter PROJ_WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_WEIGHT_PRECISION_0-1:0] mdata_out      [PROJ_WEIGHT_PARALLELISM_DIM_0 * PROJ_WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 2304;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_attention_mproj_weight [PROJ_WEIGHT_PARALLELISM_DIM_0*PROJ_WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_attention_eproj_weight;
logic folded_blocks_0_stream_blocks_11_attention_proj_weight_valid, folded_blocks_0_stream_blocks_11_attention_proj_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_attention_proj_weight_source #(
    .PROJ_WEIGHT_PRECISION_0(PROJ_WEIGHT_PRECISION_0),
    .PROJ_WEIGHT_PRECISION_1(PROJ_WEIGHT_PRECISION_1),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_0(PROJ_WEIGHT_TENSOR_SIZE_DIM_0),
    .PROJ_WEIGHT_PARALLELISM_DIM_0(PROJ_WEIGHT_PARALLELISM_DIM_0),
    .PROJ_WEIGHT_TENSOR_SIZE_DIM_1(PROJ_WEIGHT_TENSOR_SIZE_DIM_1),
    .PROJ_WEIGHT_PARALLELISM_DIM_1(PROJ_WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_attention_proj_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_attention_mproj_weight),
    .edata_out(folded_blocks_0_stream_blocks_11_attention_eproj_weight),
    .data_out_ready(folded_blocks_0_stream_blocks_11_attention_proj_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_attention_proj_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_attention_proj_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_mproj_weight: folded_blocks_0_stream_blocks_11_attention_mproj_weight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_eproj_weight: folded_blocks_0_stream_blocks_11_attention_eproj_weight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_proj_weight_valid: folded_blocks_0_stream_blocks_11_attention_proj_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_attention_proj_bias_source #(
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter PROJ_BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter PROJ_BIAS_PRECISION_0 = -1,
    parameter PROJ_BIAS_PRECISION_1 = -1,

    parameter PROJ_BIAS_PARALLELISM_DIM_0 = -1,
    parameter PROJ_BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [PROJ_BIAS_PRECISION_0-1:0] mdata_out      [PROJ_BIAS_PARALLELISM_DIM_0 * PROJ_BIAS_PARALLELISM_DIM_1-1:0],
    output logic [PROJ_BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [PROJ_BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_attention_mproj_bias [PROJ_BIAS_PARALLELISM_DIM_0*PROJ_BIAS_PARALLELISM_DIM_1 - 1:0];
logic [PROJ_BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_attention_eproj_bias;
logic folded_blocks_0_stream_blocks_11_attention_proj_bias_valid, folded_blocks_0_stream_blocks_11_attention_proj_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_attention_proj_bias_source #(
    .PROJ_BIAS_PRECISION_0(PROJ_BIAS_PRECISION_0),
    .PROJ_BIAS_PRECISION_1(PROJ_BIAS_PRECISION_1),
    .PROJ_BIAS_TENSOR_SIZE_DIM_0(PROJ_BIAS_TENSOR_SIZE_DIM_0),
    .PROJ_BIAS_PARALLELISM_DIM_0(PROJ_BIAS_PARALLELISM_DIM_0),
    .PROJ_BIAS_TENSOR_SIZE_DIM_1(PROJ_BIAS_TENSOR_SIZE_DIM_1),
    .PROJ_BIAS_PARALLELISM_DIM_1(PROJ_BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_attention_proj_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_attention_mproj_bias),
    .edata_out(folded_blocks_0_stream_blocks_11_attention_eproj_bias),
    .data_out_ready(folded_blocks_0_stream_blocks_11_attention_proj_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_attention_proj_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_attention_proj_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_mproj_bias: folded_blocks_0_stream_blocks_11_attention_mproj_bias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_eproj_bias: folded_blocks_0_stream_blocks_11_attention_eproj_bias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_attention_proj_bias_valid: folded_blocks_0_stream_blocks_11_attention_proj_bias_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_norm2_weight_source #(
    parameter WEIGHT_TENSOR_SIZE_DIM_0  = -1,
    parameter WEIGHT_TENSOR_SIZE_DIM_1  = -1,
    parameter WEIGHT_PRECISION_0 = -1,
    parameter WEIGHT_PRECISION_1 = -1,

    parameter WEIGHT_PARALLELISM_DIM_0 = -1,
    parameter WEIGHT_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [WEIGHT_PRECISION_0-1:0] mdata_out      [WEIGHT_PARALLELISM_DIM_0 * WEIGHT_PARALLELISM_DIM_1-1:0],
    output logic [WEIGHT_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [WEIGHT_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_norm2_mweight [WEIGHT_PARALLELISM_DIM_0*WEIGHT_PARALLELISM_DIM_1 - 1:0];
logic [WEIGHT_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_norm2_eweight;
logic folded_blocks_0_stream_blocks_11_norm2_weight_valid, folded_blocks_0_stream_blocks_11_norm2_weight_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_norm2_weight_source #(
    .WEIGHT_PRECISION_0(WEIGHT_PRECISION_0),
    .WEIGHT_PRECISION_1(WEIGHT_PRECISION_1),
    .WEIGHT_TENSOR_SIZE_DIM_0(WEIGHT_TENSOR_SIZE_DIM_0),
    .WEIGHT_PARALLELISM_DIM_0(WEIGHT_PARALLELISM_DIM_0),
    .WEIGHT_TENSOR_SIZE_DIM_1(WEIGHT_TENSOR_SIZE_DIM_1),
    .WEIGHT_PARALLELISM_DIM_1(WEIGHT_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_norm2_weight_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_norm2_mweight),
    .edata_out(folded_blocks_0_stream_blocks_11_norm2_eweight),
    .data_out_ready(folded_blocks_0_stream_blocks_11_norm2_weight_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_norm2_weight_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_norm2_weight_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm2_mweight: folded_blocks_0_stream_blocks_11_norm2_mweight;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm2_eweight: folded_blocks_0_stream_blocks_11_norm2_eweight;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm2_weight_valid: folded_blocks_0_stream_blocks_11_norm2_weight_valid;
end 


endmodule
        
`timescale 1ns / 1ps
module stream_blocks_11_norm2_bias_source #(
    parameter BIAS_TENSOR_SIZE_DIM_0  = -1,
    parameter BIAS_TENSOR_SIZE_DIM_1  = -1,
    parameter BIAS_PRECISION_0 = -1,
    parameter BIAS_PRECISION_1 = -1,

    parameter BIAS_PARALLELISM_DIM_0 = -1,
    parameter BIAS_PARALLELISM_DIM_1 = -1
) (
    input clk,
    input rst,

    output logic [BIAS_PRECISION_0-1:0] mdata_out      [BIAS_PARALLELISM_DIM_0 * BIAS_PARALLELISM_DIM_1-1:0],
    output logic [BIAS_PRECISION_1-1:0] edata_out,
    output logic                 data_out_valid,
    input                        data_out_ready
);
localparam REPEAT_TIMES = 1;
localparam IMAGE_DEPTH = 48;
localparam COUNTER_DEPTH = REPEAT_TIMES*IMAGE_DEPTH;
logic [$clog2(COUNTER_DEPTH) - 1 : 0] counter;

logic [BIAS_PRECISION_0 - 1:0] folded_blocks_0_stream_blocks_11_norm2_mbias [BIAS_PARALLELISM_DIM_0*BIAS_PARALLELISM_DIM_1 - 1:0];
logic [BIAS_PRECISION_1 - 1:0] folded_blocks_0_stream_blocks_11_norm2_ebias;
logic folded_blocks_0_stream_blocks_11_norm2_bias_valid, folded_blocks_0_stream_blocks_11_norm2_bias_ready;

always_ff @(posedge clk)
    if (rst) counter <= 0;
    else
        if (counter == COUNTER_DEPTH) counter <= 0;
        else if (data_out_valid && data_out_ready) counter <= counter + 1;


folded_blocks_0_stream_blocks_11_norm2_bias_source #(
    .BIAS_PRECISION_0(BIAS_PRECISION_0),
    .BIAS_PRECISION_1(BIAS_PRECISION_1),
    .BIAS_TENSOR_SIZE_DIM_0(BIAS_TENSOR_SIZE_DIM_0),
    .BIAS_PARALLELISM_DIM_0(BIAS_PARALLELISM_DIM_0),
    .BIAS_TENSOR_SIZE_DIM_1(BIAS_TENSOR_SIZE_DIM_1),
    .BIAS_PARALLELISM_DIM_1(BIAS_PARALLELISM_DIM_1)
) folded_blocks_0_stream_blocks_11_norm2_bias_source_0 (
    .clk(clk),
    .rst(rst),
    .mdata_out(folded_blocks_0_stream_blocks_11_norm2_mbias),
    .edata_out(folded_blocks_0_stream_blocks_11_norm2_ebias),
    .data_out_ready(folded_blocks_0_stream_blocks_11_norm2_bias_ready),
    .data_out_valid(folded_blocks_0_stream_blocks_11_norm2_bias_valid)
);

    


always_comb begin
    
folded_blocks_0_stream_blocks_11_norm2_bias_ready = ((0*IMAGE_DEPTH<=counter) && (counter<1*IMAGE_DEPTH))? data_out_ready:0; 
end
    
always_comb begin
    mdata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm2_mbias: folded_blocks_0_stream_blocks_11_norm2_mbias;

    edata_out = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm2_ebias: folded_blocks_0_stream_blocks_11_norm2_ebias;

    data_out_valid = (counter<IMAGE_DEPTH)?
    folded_blocks_0_stream_blocks_11_norm2_bias_valid: folded_blocks_0_stream_blocks_11_norm2_bias_valid;
end 


endmodule
        
    