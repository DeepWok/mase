
`timescale 1ns / 1ps
/* verilator lint_off UNUSEDPARAM */
module isqrt_lut #(
    parameter DATA_IN_0_PRECISION_0  = 9,
    parameter DATA_IN_0_PRECISION_1  = 7,
    parameter DATA_OUT_0_PRECISION_0 = 8,
    parameter DATA_OUT_0_PRECISION_1 = 4
) (
    /* verilator lint_off UNUSEDSIGNAL */
    input  logic [8:0] data_in_0,
    output logic [7:0] data_out_0
);


  always_comb begin
    case (data_in_0)
      9'b000000000: data_out_0 = 8'b01111111;
      9'b000000001: data_out_0 = 8'b01111111;
      9'b000000010: data_out_0 = 8'b01111111;
      9'b000000011: data_out_0 = 8'b01101000;
      9'b000000100: data_out_0 = 8'b01011010;
      9'b000000101: data_out_0 = 8'b01010001;
      9'b000000110: data_out_0 = 8'b01001010;
      9'b000000111: data_out_0 = 8'b01000100;
      9'b000001000: data_out_0 = 8'b01000000;
      9'b000001001: data_out_0 = 8'b00111100;
      9'b000001010: data_out_0 = 8'b00111001;
      9'b000001011: data_out_0 = 8'b00110111;
      9'b000001100: data_out_0 = 8'b00110100;
      9'b000001101: data_out_0 = 8'b00110010;
      9'b000001110: data_out_0 = 8'b00110000;
      9'b000001111: data_out_0 = 8'b00101111;
      9'b000010000: data_out_0 = 8'b00101101;
      9'b000010001: data_out_0 = 8'b00101100;
      9'b000010010: data_out_0 = 8'b00101011;
      9'b000010011: data_out_0 = 8'b00101010;
      9'b000010100: data_out_0 = 8'b00101000;
      9'b000010101: data_out_0 = 8'b00101000;
      9'b000010110: data_out_0 = 8'b00100111;
      9'b000010111: data_out_0 = 8'b00100110;
      9'b000011000: data_out_0 = 8'b00100101;
      9'b000011001: data_out_0 = 8'b00100100;
      9'b000011010: data_out_0 = 8'b00100011;
      9'b000011011: data_out_0 = 8'b00100011;
      9'b000011100: data_out_0 = 8'b00100010;
      9'b000011101: data_out_0 = 8'b00100010;
      9'b000011110: data_out_0 = 8'b00100001;
      9'b000011111: data_out_0 = 8'b00100001;
      9'b000100000: data_out_0 = 8'b00100000;
      9'b000100001: data_out_0 = 8'b00100000;
      9'b000100010: data_out_0 = 8'b00011111;
      9'b000100011: data_out_0 = 8'b00011111;
      9'b000100100: data_out_0 = 8'b00011110;
      9'b000100101: data_out_0 = 8'b00011110;
      9'b000100110: data_out_0 = 8'b00011101;
      9'b000100111: data_out_0 = 8'b00011101;
      9'b000101000: data_out_0 = 8'b00011101;
      9'b000101001: data_out_0 = 8'b00011100;
      9'b000101010: data_out_0 = 8'b00011100;
      9'b000101011: data_out_0 = 8'b00011100;
      9'b000101100: data_out_0 = 8'b00011011;
      9'b000101101: data_out_0 = 8'b00011011;
      9'b000101110: data_out_0 = 8'b00011011;
      9'b000101111: data_out_0 = 8'b00011010;
      9'b000110000: data_out_0 = 8'b00011010;
      9'b000110001: data_out_0 = 8'b00011010;
      9'b000110010: data_out_0 = 8'b00011010;
      9'b000110011: data_out_0 = 8'b00011001;
      9'b000110100: data_out_0 = 8'b00011001;
      9'b000110101: data_out_0 = 8'b00011001;
      9'b000110110: data_out_0 = 8'b00011001;
      9'b000110111: data_out_0 = 8'b00011000;
      9'b000111000: data_out_0 = 8'b00011000;
      9'b000111001: data_out_0 = 8'b00011000;
      9'b000111010: data_out_0 = 8'b00011000;
      9'b000111011: data_out_0 = 8'b00011000;
      9'b000111100: data_out_0 = 8'b00010111;
      9'b000111101: data_out_0 = 8'b00010111;
      9'b000111110: data_out_0 = 8'b00010111;
      9'b000111111: data_out_0 = 8'b00010111;
      9'b001000000: data_out_0 = 8'b00010111;
      9'b001000001: data_out_0 = 8'b00010110;
      9'b001000010: data_out_0 = 8'b00010110;
      9'b001000011: data_out_0 = 8'b00010110;
      9'b001000100: data_out_0 = 8'b00010110;
      9'b001000101: data_out_0 = 8'b00010110;
      9'b001000110: data_out_0 = 8'b00010110;
      9'b001000111: data_out_0 = 8'b00010101;
      9'b001001000: data_out_0 = 8'b00010101;
      9'b001001001: data_out_0 = 8'b00010101;
      9'b001001010: data_out_0 = 8'b00010101;
      9'b001001011: data_out_0 = 8'b00010101;
      9'b001001100: data_out_0 = 8'b00010101;
      9'b001001101: data_out_0 = 8'b00010101;
      9'b001001110: data_out_0 = 8'b00010100;
      9'b001001111: data_out_0 = 8'b00010100;
      9'b001010000: data_out_0 = 8'b00010100;
      9'b001010001: data_out_0 = 8'b00010100;
      9'b001010010: data_out_0 = 8'b00010100;
      9'b001010011: data_out_0 = 8'b00010100;
      9'b001010100: data_out_0 = 8'b00010100;
      9'b001010101: data_out_0 = 8'b00010100;
      9'b001010110: data_out_0 = 8'b00010100;
      9'b001010111: data_out_0 = 8'b00010011;
      9'b001011000: data_out_0 = 8'b00010011;
      9'b001011001: data_out_0 = 8'b00010011;
      9'b001011010: data_out_0 = 8'b00010011;
      9'b001011011: data_out_0 = 8'b00010011;
      9'b001011100: data_out_0 = 8'b00010011;
      9'b001011101: data_out_0 = 8'b00010011;
      9'b001011110: data_out_0 = 8'b00010011;
      9'b001011111: data_out_0 = 8'b00010011;
      9'b001100000: data_out_0 = 8'b00010010;
      9'b001100001: data_out_0 = 8'b00010010;
      9'b001100010: data_out_0 = 8'b00010010;
      9'b001100011: data_out_0 = 8'b00010010;
      9'b001100100: data_out_0 = 8'b00010010;
      9'b001100101: data_out_0 = 8'b00010010;
      9'b001100110: data_out_0 = 8'b00010010;
      9'b001100111: data_out_0 = 8'b00010010;
      9'b001101000: data_out_0 = 8'b00010010;
      9'b001101001: data_out_0 = 8'b00010010;
      9'b001101010: data_out_0 = 8'b00010010;
      9'b001101011: data_out_0 = 8'b00010001;
      9'b001101100: data_out_0 = 8'b00010001;
      9'b001101101: data_out_0 = 8'b00010001;
      9'b001101110: data_out_0 = 8'b00010001;
      9'b001101111: data_out_0 = 8'b00010001;
      9'b001110000: data_out_0 = 8'b00010001;
      9'b001110001: data_out_0 = 8'b00010001;
      9'b001110010: data_out_0 = 8'b00010001;
      9'b001110011: data_out_0 = 8'b00010001;
      9'b001110100: data_out_0 = 8'b00010001;
      9'b001110101: data_out_0 = 8'b00010001;
      9'b001110110: data_out_0 = 8'b00010001;
      9'b001110111: data_out_0 = 8'b00010001;
      9'b001111000: data_out_0 = 8'b00010001;
      9'b001111001: data_out_0 = 8'b00010000;
      9'b001111010: data_out_0 = 8'b00010000;
      9'b001111011: data_out_0 = 8'b00010000;
      9'b001111100: data_out_0 = 8'b00010000;
      9'b001111101: data_out_0 = 8'b00010000;
      9'b001111110: data_out_0 = 8'b00010000;
      9'b001111111: data_out_0 = 8'b00010000;
      9'b010000000: data_out_0 = 8'b00010000;
      9'b010000001: data_out_0 = 8'b00010000;
      9'b010000010: data_out_0 = 8'b00010000;
      9'b010000011: data_out_0 = 8'b00010000;
      9'b010000100: data_out_0 = 8'b00010000;
      9'b010000101: data_out_0 = 8'b00010000;
      9'b010000110: data_out_0 = 8'b00010000;
      9'b010000111: data_out_0 = 8'b00010000;
      9'b010001000: data_out_0 = 8'b00010000;
      9'b010001001: data_out_0 = 8'b00001111;
      9'b010001010: data_out_0 = 8'b00001111;
      9'b010001011: data_out_0 = 8'b00001111;
      9'b010001100: data_out_0 = 8'b00001111;
      9'b010001101: data_out_0 = 8'b00001111;
      9'b010001110: data_out_0 = 8'b00001111;
      9'b010001111: data_out_0 = 8'b00001111;
      9'b010010000: data_out_0 = 8'b00001111;
      9'b010010001: data_out_0 = 8'b00001111;
      9'b010010010: data_out_0 = 8'b00001111;
      9'b010010011: data_out_0 = 8'b00001111;
      9'b010010100: data_out_0 = 8'b00001111;
      9'b010010101: data_out_0 = 8'b00001111;
      9'b010010110: data_out_0 = 8'b00001111;
      9'b010010111: data_out_0 = 8'b00001111;
      9'b010011000: data_out_0 = 8'b00001111;
      9'b010011001: data_out_0 = 8'b00001111;
      9'b010011010: data_out_0 = 8'b00001111;
      9'b010011011: data_out_0 = 8'b00001111;
      9'b010011100: data_out_0 = 8'b00001110;
      9'b010011101: data_out_0 = 8'b00001110;
      9'b010011110: data_out_0 = 8'b00001110;
      9'b010011111: data_out_0 = 8'b00001110;
      9'b010100000: data_out_0 = 8'b00001110;
      9'b010100001: data_out_0 = 8'b00001110;
      9'b010100010: data_out_0 = 8'b00001110;
      9'b010100011: data_out_0 = 8'b00001110;
      9'b010100100: data_out_0 = 8'b00001110;
      9'b010100101: data_out_0 = 8'b00001110;
      9'b010100110: data_out_0 = 8'b00001110;
      9'b010100111: data_out_0 = 8'b00001110;
      9'b010101000: data_out_0 = 8'b00001110;
      9'b010101001: data_out_0 = 8'b00001110;
      9'b010101010: data_out_0 = 8'b00001110;
      9'b010101011: data_out_0 = 8'b00001110;
      9'b010101100: data_out_0 = 8'b00001110;
      9'b010101101: data_out_0 = 8'b00001110;
      9'b010101110: data_out_0 = 8'b00001110;
      9'b010101111: data_out_0 = 8'b00001110;
      9'b010110000: data_out_0 = 8'b00001110;
      9'b010110001: data_out_0 = 8'b00001110;
      9'b010110010: data_out_0 = 8'b00001110;
      9'b010110011: data_out_0 = 8'b00001110;
      9'b010110100: data_out_0 = 8'b00001101;
      9'b010110101: data_out_0 = 8'b00001101;
      9'b010110110: data_out_0 = 8'b00001101;
      9'b010110111: data_out_0 = 8'b00001101;
      9'b010111000: data_out_0 = 8'b00001101;
      9'b010111001: data_out_0 = 8'b00001101;
      9'b010111010: data_out_0 = 8'b00001101;
      9'b010111011: data_out_0 = 8'b00001101;
      9'b010111100: data_out_0 = 8'b00001101;
      9'b010111101: data_out_0 = 8'b00001101;
      9'b010111110: data_out_0 = 8'b00001101;
      9'b010111111: data_out_0 = 8'b00001101;
      9'b011000000: data_out_0 = 8'b00001101;
      9'b011000001: data_out_0 = 8'b00001101;
      9'b011000010: data_out_0 = 8'b00001101;
      9'b011000011: data_out_0 = 8'b00001101;
      9'b011000100: data_out_0 = 8'b00001101;
      9'b011000101: data_out_0 = 8'b00001101;
      9'b011000110: data_out_0 = 8'b00001101;
      9'b011000111: data_out_0 = 8'b00001101;
      9'b011001000: data_out_0 = 8'b00001101;
      9'b011001001: data_out_0 = 8'b00001101;
      9'b011001010: data_out_0 = 8'b00001101;
      9'b011001011: data_out_0 = 8'b00001101;
      9'b011001100: data_out_0 = 8'b00001101;
      9'b011001101: data_out_0 = 8'b00001101;
      9'b011001110: data_out_0 = 8'b00001101;
      9'b011001111: data_out_0 = 8'b00001101;
      9'b011010000: data_out_0 = 8'b00001101;
      9'b011010001: data_out_0 = 8'b00001101;
      9'b011010010: data_out_0 = 8'b00001100;
      9'b011010011: data_out_0 = 8'b00001100;
      9'b011010100: data_out_0 = 8'b00001100;
      9'b011010101: data_out_0 = 8'b00001100;
      9'b011010110: data_out_0 = 8'b00001100;
      9'b011010111: data_out_0 = 8'b00001100;
      9'b011011000: data_out_0 = 8'b00001100;
      9'b011011001: data_out_0 = 8'b00001100;
      9'b011011010: data_out_0 = 8'b00001100;
      9'b011011011: data_out_0 = 8'b00001100;
      9'b011011100: data_out_0 = 8'b00001100;
      9'b011011101: data_out_0 = 8'b00001100;
      9'b011011110: data_out_0 = 8'b00001100;
      9'b011011111: data_out_0 = 8'b00001100;
      9'b011100000: data_out_0 = 8'b00001100;
      9'b011100001: data_out_0 = 8'b00001100;
      9'b011100010: data_out_0 = 8'b00001100;
      9'b011100011: data_out_0 = 8'b00001100;
      9'b011100100: data_out_0 = 8'b00001100;
      9'b011100101: data_out_0 = 8'b00001100;
      9'b011100110: data_out_0 = 8'b00001100;
      9'b011100111: data_out_0 = 8'b00001100;
      9'b011101000: data_out_0 = 8'b00001100;
      9'b011101001: data_out_0 = 8'b00001100;
      9'b011101010: data_out_0 = 8'b00001100;
      9'b011101011: data_out_0 = 8'b00001100;
      9'b011101100: data_out_0 = 8'b00001100;
      9'b011101101: data_out_0 = 8'b00001100;
      9'b011101110: data_out_0 = 8'b00001100;
      9'b011101111: data_out_0 = 8'b00001100;
      9'b011110000: data_out_0 = 8'b00001100;
      9'b011110001: data_out_0 = 8'b00001100;
      9'b011110010: data_out_0 = 8'b00001100;
      9'b011110011: data_out_0 = 8'b00001100;
      9'b011110100: data_out_0 = 8'b00001100;
      9'b011110101: data_out_0 = 8'b00001100;
      9'b011110110: data_out_0 = 8'b00001100;
      9'b011110111: data_out_0 = 8'b00001100;
      9'b011111000: data_out_0 = 8'b00001011;
      9'b011111001: data_out_0 = 8'b00001011;
      9'b011111010: data_out_0 = 8'b00001011;
      9'b011111011: data_out_0 = 8'b00001011;
      9'b011111100: data_out_0 = 8'b00001011;
      9'b011111101: data_out_0 = 8'b00001011;
      9'b011111110: data_out_0 = 8'b00001011;
      9'b011111111: data_out_0 = 8'b00001011;
      default: data_out_0 = 8'b0;
    endcase
  end
endmodule
